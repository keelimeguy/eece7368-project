-- Keelin Becker-Wheeler
-- lut_square_ticks.vhd

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity lut_square_ticks is
    port (
        freq              : in  std_logic_vector(13 downto 0);
        half_period_ticks : out integer
    );
end lut_square_ticks;

architecture Behavioral of lut_square_ticks is
begin
    with freq select
        half_period_ticks <= 0 when "00000000000000",
                             50000000 when "00000000000001",
                             25000000 when "00000000000010",
                             16666667 when "00000000000011",
                             12500000 when "00000000000100",
                             10000000 when "00000000000101",
                             8333333 when "00000000000110",
                             7142857 when "00000000000111",
                             6250000 when "00000000001000",
                             5555556 when "00000000001001",
                             5000000 when "00000000001010",
                             4545455 when "00000000001011",
                             4166667 when "00000000001100",
                             3846154 when "00000000001101",
                             3571429 when "00000000001110",
                             3333333 when "00000000001111",
                             3125000 when "00000000010000",
                             2941176 when "00000000010001",
                             2777778 when "00000000010010",
                             2631579 when "00000000010011",
                             2500000 when "00000000010100",
                             2380952 when "00000000010101",
                             2272727 when "00000000010110",
                             2173913 when "00000000010111",
                             2083333 when "00000000011000",
                             2000000 when "00000000011001",
                             1923077 when "00000000011010",
                             1851852 when "00000000011011",
                             1785714 when "00000000011100",
                             1724138 when "00000000011101",
                             1666667 when "00000000011110",
                             1612903 when "00000000011111",
                             1562500 when "00000000100000",
                             1515152 when "00000000100001",
                             1470588 when "00000000100010",
                             1428571 when "00000000100011",
                             1388889 when "00000000100100",
                             1351351 when "00000000100101",
                             1315789 when "00000000100110",
                             1282051 when "00000000100111",
                             1250000 when "00000000101000",
                             1219512 when "00000000101001",
                             1190476 when "00000000101010",
                             1162791 when "00000000101011",
                             1136364 when "00000000101100",
                             1111111 when "00000000101101",
                             1086957 when "00000000101110",
                             1063830 when "00000000101111",
                             1041667 when "00000000110000",
                             1020408 when "00000000110001",
                             1000000 when "00000000110010",
                             980392 when "00000000110011",
                             961538 when "00000000110100",
                             943396 when "00000000110101",
                             925926 when "00000000110110",
                             909091 when "00000000110111",
                             892857 when "00000000111000",
                             877193 when "00000000111001",
                             862069 when "00000000111010",
                             847458 when "00000000111011",
                             833333 when "00000000111100",
                             819672 when "00000000111101",
                             806452 when "00000000111110",
                             793651 when "00000000111111",
                             781250 when "00000001000000",
                             769231 when "00000001000001",
                             757576 when "00000001000010",
                             746269 when "00000001000011",
                             735294 when "00000001000100",
                             724638 when "00000001000101",
                             714286 when "00000001000110",
                             704225 when "00000001000111",
                             694444 when "00000001001000",
                             684932 when "00000001001001",
                             675676 when "00000001001010",
                             666667 when "00000001001011",
                             657895 when "00000001001100",
                             649351 when "00000001001101",
                             641026 when "00000001001110",
                             632911 when "00000001001111",
                             625000 when "00000001010000",
                             617284 when "00000001010001",
                             609756 when "00000001010010",
                             602410 when "00000001010011",
                             595238 when "00000001010100",
                             588235 when "00000001010101",
                             581395 when "00000001010110",
                             574713 when "00000001010111",
                             568182 when "00000001011000",
                             561798 when "00000001011001",
                             555556 when "00000001011010",
                             549451 when "00000001011011",
                             543478 when "00000001011100",
                             537634 when "00000001011101",
                             531915 when "00000001011110",
                             526316 when "00000001011111",
                             520833 when "00000001100000",
                             515464 when "00000001100001",
                             510204 when "00000001100010",
                             505051 when "00000001100011",
                             500000 when "00000001100100",
                             495050 when "00000001100101",
                             490196 when "00000001100110",
                             485437 when "00000001100111",
                             480769 when "00000001101000",
                             476190 when "00000001101001",
                             471698 when "00000001101010",
                             467290 when "00000001101011",
                             462963 when "00000001101100",
                             458716 when "00000001101101",
                             454545 when "00000001101110",
                             450450 when "00000001101111",
                             446429 when "00000001110000",
                             442478 when "00000001110001",
                             438596 when "00000001110010",
                             434783 when "00000001110011",
                             431034 when "00000001110100",
                             427350 when "00000001110101",
                             423729 when "00000001110110",
                             420168 when "00000001110111",
                             416667 when "00000001111000",
                             413223 when "00000001111001",
                             409836 when "00000001111010",
                             406504 when "00000001111011",
                             403226 when "00000001111100",
                             400000 when "00000001111101",
                             396825 when "00000001111110",
                             393701 when "00000001111111",
                             390625 when "00000010000000",
                             387597 when "00000010000001",
                             384615 when "00000010000010",
                             381679 when "00000010000011",
                             378788 when "00000010000100",
                             375940 when "00000010000101",
                             373134 when "00000010000110",
                             370370 when "00000010000111",
                             367647 when "00000010001000",
                             364964 when "00000010001001",
                             362319 when "00000010001010",
                             359712 when "00000010001011",
                             357143 when "00000010001100",
                             354610 when "00000010001101",
                             352113 when "00000010001110",
                             349650 when "00000010001111",
                             347222 when "00000010010000",
                             344828 when "00000010010001",
                             342466 when "00000010010010",
                             340136 when "00000010010011",
                             337838 when "00000010010100",
                             335570 when "00000010010101",
                             333333 when "00000010010110",
                             331126 when "00000010010111",
                             328947 when "00000010011000",
                             326797 when "00000010011001",
                             324675 when "00000010011010",
                             322581 when "00000010011011",
                             320513 when "00000010011100",
                             318471 when "00000010011101",
                             316456 when "00000010011110",
                             314465 when "00000010011111",
                             312500 when "00000010100000",
                             310559 when "00000010100001",
                             308642 when "00000010100010",
                             306748 when "00000010100011",
                             304878 when "00000010100100",
                             303030 when "00000010100101",
                             301205 when "00000010100110",
                             299401 when "00000010100111",
                             297619 when "00000010101000",
                             295858 when "00000010101001",
                             294118 when "00000010101010",
                             292398 when "00000010101011",
                             290698 when "00000010101100",
                             289017 when "00000010101101",
                             287356 when "00000010101110",
                             285714 when "00000010101111",
                             284091 when "00000010110000",
                             282486 when "00000010110001",
                             280899 when "00000010110010",
                             279330 when "00000010110011",
                             277778 when "00000010110100",
                             276243 when "00000010110101",
                             274725 when "00000010110110",
                             273224 when "00000010110111",
                             271739 when "00000010111000",
                             270270 when "00000010111001",
                             268817 when "00000010111010",
                             267380 when "00000010111011",
                             265957 when "00000010111100",
                             264550 when "00000010111101",
                             263158 when "00000010111110",
                             261780 when "00000010111111",
                             260417 when "00000011000000",
                             259067 when "00000011000001",
                             257732 when "00000011000010",
                             256410 when "00000011000011",
                             255102 when "00000011000100",
                             253807 when "00000011000101",
                             252525 when "00000011000110",
                             251256 when "00000011000111",
                             250000 when "00000011001000",
                             248756 when "00000011001001",
                             247525 when "00000011001010",
                             246305 when "00000011001011",
                             245098 when "00000011001100",
                             243902 when "00000011001101",
                             242718 when "00000011001110",
                             241546 when "00000011001111",
                             240385 when "00000011010000",
                             239234 when "00000011010001",
                             238095 when "00000011010010",
                             236967 when "00000011010011",
                             235849 when "00000011010100",
                             234742 when "00000011010101",
                             233645 when "00000011010110",
                             232558 when "00000011010111",
                             231481 when "00000011011000",
                             230415 when "00000011011001",
                             229358 when "00000011011010",
                             228311 when "00000011011011",
                             227273 when "00000011011100",
                             226244 when "00000011011101",
                             225225 when "00000011011110",
                             224215 when "00000011011111",
                             223214 when "00000011100000",
                             222222 when "00000011100001",
                             221239 when "00000011100010",
                             220264 when "00000011100011",
                             219298 when "00000011100100",
                             218341 when "00000011100101",
                             217391 when "00000011100110",
                             216450 when "00000011100111",
                             215517 when "00000011101000",
                             214592 when "00000011101001",
                             213675 when "00000011101010",
                             212766 when "00000011101011",
                             211864 when "00000011101100",
                             210970 when "00000011101101",
                             210084 when "00000011101110",
                             209205 when "00000011101111",
                             208333 when "00000011110000",
                             207469 when "00000011110001",
                             206612 when "00000011110010",
                             205761 when "00000011110011",
                             204918 when "00000011110100",
                             204082 when "00000011110101",
                             203252 when "00000011110110",
                             202429 when "00000011110111",
                             201613 when "00000011111000",
                             200803 when "00000011111001",
                             200000 when "00000011111010",
                             199203 when "00000011111011",
                             198413 when "00000011111100",
                             197628 when "00000011111101",
                             196850 when "00000011111110",
                             196078 when "00000011111111",
                             195313 when "00000100000000",
                             194553 when "00000100000001",
                             193798 when "00000100000010",
                             193050 when "00000100000011",
                             192308 when "00000100000100",
                             191571 when "00000100000101",
                             190840 when "00000100000110",
                             190114 when "00000100000111",
                             189394 when "00000100001000",
                             188679 when "00000100001001",
                             187970 when "00000100001010",
                             187266 when "00000100001011",
                             186567 when "00000100001100",
                             185874 when "00000100001101",
                             185185 when "00000100001110",
                             184502 when "00000100001111",
                             183824 when "00000100010000",
                             183150 when "00000100010001",
                             182482 when "00000100010010",
                             181818 when "00000100010011",
                             181159 when "00000100010100",
                             180505 when "00000100010101",
                             179856 when "00000100010110",
                             179211 when "00000100010111",
                             178571 when "00000100011000",
                             177936 when "00000100011001",
                             177305 when "00000100011010",
                             176678 when "00000100011011",
                             176056 when "00000100011100",
                             175439 when "00000100011101",
                             174825 when "00000100011110",
                             174216 when "00000100011111",
                             173611 when "00000100100000",
                             173010 when "00000100100001",
                             172414 when "00000100100010",
                             171821 when "00000100100011",
                             171233 when "00000100100100",
                             170648 when "00000100100101",
                             170068 when "00000100100110",
                             169492 when "00000100100111",
                             168919 when "00000100101000",
                             168350 when "00000100101001",
                             167785 when "00000100101010",
                             167224 when "00000100101011",
                             166667 when "00000100101100",
                             166113 when "00000100101101",
                             165563 when "00000100101110",
                             165017 when "00000100101111",
                             164474 when "00000100110000",
                             163934 when "00000100110001",
                             163399 when "00000100110010",
                             162866 when "00000100110011",
                             162338 when "00000100110100",
                             161812 when "00000100110101",
                             161290 when "00000100110110",
                             160772 when "00000100110111",
                             160256 when "00000100111000",
                             159744 when "00000100111001",
                             159236 when "00000100111010",
                             158730 when "00000100111011",
                             158228 when "00000100111100",
                             157729 when "00000100111101",
                             157233 when "00000100111110",
                             156740 when "00000100111111",
                             156250 when "00000101000000",
                             155763 when "00000101000001",
                             155280 when "00000101000010",
                             154799 when "00000101000011",
                             154321 when "00000101000100",
                             153846 when "00000101000101",
                             153374 when "00000101000110",
                             152905 when "00000101000111",
                             152439 when "00000101001000",
                             151976 when "00000101001001",
                             151515 when "00000101001010",
                             151057 when "00000101001011",
                             150602 when "00000101001100",
                             150150 when "00000101001101",
                             149701 when "00000101001110",
                             149254 when "00000101001111",
                             148810 when "00000101010000",
                             148368 when "00000101010001",
                             147929 when "00000101010010",
                             147493 when "00000101010011",
                             147059 when "00000101010100",
                             146628 when "00000101010101",
                             146199 when "00000101010110",
                             145773 when "00000101010111",
                             145349 when "00000101011000",
                             144928 when "00000101011001",
                             144509 when "00000101011010",
                             144092 when "00000101011011",
                             143678 when "00000101011100",
                             143266 when "00000101011101",
                             142857 when "00000101011110",
                             142450 when "00000101011111",
                             142045 when "00000101100000",
                             141643 when "00000101100001",
                             141243 when "00000101100010",
                             140845 when "00000101100011",
                             140449 when "00000101100100",
                             140056 when "00000101100101",
                             139665 when "00000101100110",
                             139276 when "00000101100111",
                             138889 when "00000101101000",
                             138504 when "00000101101001",
                             138122 when "00000101101010",
                             137741 when "00000101101011",
                             137363 when "00000101101100",
                             136986 when "00000101101101",
                             136612 when "00000101101110",
                             136240 when "00000101101111",
                             135870 when "00000101110000",
                             135501 when "00000101110001",
                             135135 when "00000101110010",
                             134771 when "00000101110011",
                             134409 when "00000101110100",
                             134048 when "00000101110101",
                             133690 when "00000101110110",
                             133333 when "00000101110111",
                             132979 when "00000101111000",
                             132626 when "00000101111001",
                             132275 when "00000101111010",
                             131926 when "00000101111011",
                             131579 when "00000101111100",
                             131234 when "00000101111101",
                             130890 when "00000101111110",
                             130548 when "00000101111111",
                             130208 when "00000110000000",
                             129870 when "00000110000001",
                             129534 when "00000110000010",
                             129199 when "00000110000011",
                             128866 when "00000110000100",
                             128535 when "00000110000101",
                             128205 when "00000110000110",
                             127877 when "00000110000111",
                             127551 when "00000110001000",
                             127226 when "00000110001001",
                             126904 when "00000110001010",
                             126582 when "00000110001011",
                             126263 when "00000110001100",
                             125945 when "00000110001101",
                             125628 when "00000110001110",
                             125313 when "00000110001111",
                             125000 when "00000110010000",
                             124688 when "00000110010001",
                             124378 when "00000110010010",
                             124069 when "00000110010011",
                             123762 when "00000110010100",
                             123457 when "00000110010101",
                             123153 when "00000110010110",
                             122850 when "00000110010111",
                             122549 when "00000110011000",
                             122249 when "00000110011001",
                             121951 when "00000110011010",
                             121655 when "00000110011011",
                             121359 when "00000110011100",
                             121065 when "00000110011101",
                             120773 when "00000110011110",
                             120482 when "00000110011111",
                             120192 when "00000110100000",
                             119904 when "00000110100001",
                             119617 when "00000110100010",
                             119332 when "00000110100011",
                             119048 when "00000110100100",
                             118765 when "00000110100101",
                             118483 when "00000110100110",
                             118203 when "00000110100111",
                             117925 when "00000110101000",
                             117647 when "00000110101001",
                             117371 when "00000110101010",
                             117096 when "00000110101011",
                             116822 when "00000110101100",
                             116550 when "00000110101101",
                             116279 when "00000110101110",
                             116009 when "00000110101111",
                             115741 when "00000110110000",
                             115473 when "00000110110001",
                             115207 when "00000110110010",
                             114943 when "00000110110011",
                             114679 when "00000110110100",
                             114416 when "00000110110101",
                             114155 when "00000110110110",
                             113895 when "00000110110111",
                             113636 when "00000110111000",
                             113379 when "00000110111001",
                             113122 when "00000110111010",
                             112867 when "00000110111011",
                             112613 when "00000110111100",
                             112360 when "00000110111101",
                             112108 when "00000110111110",
                             111857 when "00000110111111",
                             111607 when "00000111000000",
                             111359 when "00000111000001",
                             111111 when "00000111000010",
                             110865 when "00000111000011",
                             110619 when "00000111000100",
                             110375 when "00000111000101",
                             110132 when "00000111000110",
                             109890 when "00000111000111",
                             109649 when "00000111001000",
                             109409 when "00000111001001",
                             109170 when "00000111001010",
                             108932 when "00000111001011",
                             108696 when "00000111001100",
                             108460 when "00000111001101",
                             108225 when "00000111001110",
                             107991 when "00000111001111",
                             107759 when "00000111010000",
                             107527 when "00000111010001",
                             107296 when "00000111010010",
                             107066 when "00000111010011",
                             106838 when "00000111010100",
                             106610 when "00000111010101",
                             106383 when "00000111010110",
                             106157 when "00000111010111",
                             105932 when "00000111011000",
                             105708 when "00000111011001",
                             105485 when "00000111011010",
                             105263 when "00000111011011",
                             105042 when "00000111011100",
                             104822 when "00000111011101",
                             104603 when "00000111011110",
                             104384 when "00000111011111",
                             104167 when "00000111100000",
                             103950 when "00000111100001",
                             103734 when "00000111100010",
                             103520 when "00000111100011",
                             103306 when "00000111100100",
                             103093 when "00000111100101",
                             102881 when "00000111100110",
                             102669 when "00000111100111",
                             102459 when "00000111101000",
                             102249 when "00000111101001",
                             102041 when "00000111101010",
                             101833 when "00000111101011",
                             101626 when "00000111101100",
                             101420 when "00000111101101",
                             101215 when "00000111101110",
                             101010 when "00000111101111",
                             100806 when "00000111110000",
                             100604 when "00000111110001",
                             100402 when "00000111110010",
                             100200 when "00000111110011",
                             100000 when "00000111110100",
                             99800 when "00000111110101",
                             99602 when "00000111110110",
                             99404 when "00000111110111",
                             99206 when "00000111111000",
                             99010 when "00000111111001",
                             98814 when "00000111111010",
                             98619 when "00000111111011",
                             98425 when "00000111111100",
                             98232 when "00000111111101",
                             98039 when "00000111111110",
                             97847 when "00000111111111",
                             97656 when "00001000000000",
                             97466 when "00001000000001",
                             97276 when "00001000000010",
                             97087 when "00001000000011",
                             96899 when "00001000000100",
                             96712 when "00001000000101",
                             96525 when "00001000000110",
                             96339 when "00001000000111",
                             96154 when "00001000001000",
                             95969 when "00001000001001",
                             95785 when "00001000001010",
                             95602 when "00001000001011",
                             95420 when "00001000001100",
                             95238 when "00001000001101",
                             95057 when "00001000001110",
                             94877 when "00001000001111",
                             94697 when "00001000010000",
                             94518 when "00001000010001",
                             94340 when "00001000010010",
                             94162 when "00001000010011",
                             93985 when "00001000010100",
                             93809 when "00001000010101",
                             93633 when "00001000010110",
                             93458 when "00001000010111",
                             93284 when "00001000011000",
                             93110 when "00001000011001",
                             92937 when "00001000011010",
                             92764 when "00001000011011",
                             92593 when "00001000011100",
                             92421 when "00001000011101",
                             92251 when "00001000011110",
                             92081 when "00001000011111",
                             91912 when "00001000100000",
                             91743 when "00001000100001",
                             91575 when "00001000100010",
                             91408 when "00001000100011",
                             91241 when "00001000100100",
                             91075 when "00001000100101",
                             90909 when "00001000100110",
                             90744 when "00001000100111",
                             90580 when "00001000101000",
                             90416 when "00001000101001",
                             90253 when "00001000101010",
                             90090 when "00001000101011",
                             89928 when "00001000101100",
                             89767 when "00001000101101",
                             89606 when "00001000101110",
                             89445 when "00001000101111",
                             89286 when "00001000110000",
                             89127 when "00001000110001",
                             88968 when "00001000110010",
                             88810 when "00001000110011",
                             88652 when "00001000110100",
                             88496 when "00001000110101",
                             88339 when "00001000110110",
                             88183 when "00001000110111",
                             88028 when "00001000111000",
                             87873 when "00001000111001",
                             87719 when "00001000111010",
                             87566 when "00001000111011",
                             87413 when "00001000111100",
                             87260 when "00001000111101",
                             87108 when "00001000111110",
                             86957 when "00001000111111",
                             86806 when "00001001000000",
                             86655 when "00001001000001",
                             86505 when "00001001000010",
                             86356 when "00001001000011",
                             86207 when "00001001000100",
                             86059 when "00001001000101",
                             85911 when "00001001000110",
                             85763 when "00001001000111",
                             85616 when "00001001001000",
                             85470 when "00001001001001",
                             85324 when "00001001001010",
                             85179 when "00001001001011",
                             85034 when "00001001001100",
                             84890 when "00001001001101",
                             84746 when "00001001001110",
                             84602 when "00001001001111",
                             84459 when "00001001010000",
                             84317 when "00001001010001",
                             84175 when "00001001010010",
                             84034 when "00001001010011",
                             83893 when "00001001010100",
                             83752 when "00001001010101",
                             83612 when "00001001010110",
                             83472 when "00001001010111",
                             83333 when "00001001011000",
                             83195 when "00001001011001",
                             83056 when "00001001011010",
                             82919 when "00001001011011",
                             82781 when "00001001011100",
                             82645 when "00001001011101",
                             82508 when "00001001011110",
                             82372 when "00001001011111",
                             82237 when "00001001100000",
                             82102 when "00001001100001",
                             81967 when "00001001100010",
                             81833 when "00001001100011",
                             81699 when "00001001100100",
                             81566 when "00001001100101",
                             81433 when "00001001100110",
                             81301 when "00001001100111",
                             81169 when "00001001101000",
                             81037 when "00001001101001",
                             80906 when "00001001101010",
                             80775 when "00001001101011",
                             80645 when "00001001101100",
                             80515 when "00001001101101",
                             80386 when "00001001101110",
                             80257 when "00001001101111",
                             80128 when "00001001110000",
                             80000 when "00001001110001",
                             79872 when "00001001110010",
                             79745 when "00001001110011",
                             79618 when "00001001110100",
                             79491 when "00001001110101",
                             79365 when "00001001110110",
                             79239 when "00001001110111",
                             79114 when "00001001111000",
                             78989 when "00001001111001",
                             78864 when "00001001111010",
                             78740 when "00001001111011",
                             78616 when "00001001111100",
                             78493 when "00001001111101",
                             78370 when "00001001111110",
                             78247 when "00001001111111",
                             78125 when "00001010000000",
                             78003 when "00001010000001",
                             77882 when "00001010000010",
                             77760 when "00001010000011",
                             77640 when "00001010000100",
                             77519 when "00001010000101",
                             77399 when "00001010000110",
                             77280 when "00001010000111",
                             77160 when "00001010001000",
                             77042 when "00001010001001",
                             76923 when "00001010001010",
                             76805 when "00001010001011",
                             76687 when "00001010001100",
                             76570 when "00001010001101",
                             76453 when "00001010001110",
                             76336 when "00001010001111",
                             76220 when "00001010010000",
                             76104 when "00001010010001",
                             75988 when "00001010010010",
                             75873 when "00001010010011",
                             75758 when "00001010010100",
                             75643 when "00001010010101",
                             75529 when "00001010010110",
                             75415 when "00001010010111",
                             75301 when "00001010011000",
                             75188 when "00001010011001",
                             75075 when "00001010011010",
                             74963 when "00001010011011",
                             74850 when "00001010011100",
                             74738 when "00001010011101",
                             74627 when "00001010011110",
                             74516 when "00001010011111",
                             74405 when "00001010100000",
                             74294 when "00001010100001",
                             74184 when "00001010100010",
                             74074 when "00001010100011",
                             73964 when "00001010100100",
                             73855 when "00001010100101",
                             73746 when "00001010100110",
                             73638 when "00001010100111",
                             73529 when "00001010101000",
                             73421 when "00001010101001",
                             73314 when "00001010101010",
                             73206 when "00001010101011",
                             73099 when "00001010101100",
                             72993 when "00001010101101",
                             72886 when "00001010101110",
                             72780 when "00001010101111",
                             72674 when "00001010110000",
                             72569 when "00001010110001",
                             72464 when "00001010110010",
                             72359 when "00001010110011",
                             72254 when "00001010110100",
                             72150 when "00001010110101",
                             72046 when "00001010110110",
                             71942 when "00001010110111",
                             71839 when "00001010111000",
                             71736 when "00001010111001",
                             71633 when "00001010111010",
                             71531 when "00001010111011",
                             71429 when "00001010111100",
                             71327 when "00001010111101",
                             71225 when "00001010111110",
                             71124 when "00001010111111",
                             71023 when "00001011000000",
                             70922 when "00001011000001",
                             70822 when "00001011000010",
                             70721 when "00001011000011",
                             70621 when "00001011000100",
                             70522 when "00001011000101",
                             70423 when "00001011000110",
                             70323 when "00001011000111",
                             70225 when "00001011001000",
                             70126 when "00001011001001",
                             70028 when "00001011001010",
                             69930 when "00001011001011",
                             69832 when "00001011001100",
                             69735 when "00001011001101",
                             69638 when "00001011001110",
                             69541 when "00001011001111",
                             69444 when "00001011010000",
                             69348 when "00001011010001",
                             69252 when "00001011010010",
                             69156 when "00001011010011",
                             69061 when "00001011010100",
                             68966 when "00001011010101",
                             68871 when "00001011010110",
                             68776 when "00001011010111",
                             68681 when "00001011011000",
                             68587 when "00001011011001",
                             68493 when "00001011011010",
                             68399 when "00001011011011",
                             68306 when "00001011011100",
                             68213 when "00001011011101",
                             68120 when "00001011011110",
                             68027 when "00001011011111",
                             67935 when "00001011100000",
                             67843 when "00001011100001",
                             67751 when "00001011100010",
                             67659 when "00001011100011",
                             67568 when "00001011100100",
                             67476 when "00001011100101",
                             67385 when "00001011100110",
                             67295 when "00001011100111",
                             67204 when "00001011101000",
                             67114 when "00001011101001",
                             67024 when "00001011101010",
                             66934 when "00001011101011",
                             66845 when "00001011101100",
                             66756 when "00001011101101",
                             66667 when "00001011101110",
                             66578 when "00001011101111",
                             66489 when "00001011110000",
                             66401 when "00001011110001",
                             66313 when "00001011110010",
                             66225 when "00001011110011",
                             66138 when "00001011110100",
                             66050 when "00001011110101",
                             65963 when "00001011110110",
                             65876 when "00001011110111",
                             65789 when "00001011111000",
                             65703 when "00001011111001",
                             65617 when "00001011111010",
                             65531 when "00001011111011",
                             65445 when "00001011111100",
                             65359 when "00001011111101",
                             65274 when "00001011111110",
                             65189 when "00001011111111",
                             65104 when "00001100000000",
                             65020 when "00001100000001",
                             64935 when "00001100000010",
                             64851 when "00001100000011",
                             64767 when "00001100000100",
                             64683 when "00001100000101",
                             64599 when "00001100000110",
                             64516 when "00001100000111",
                             64433 when "00001100001000",
                             64350 when "00001100001001",
                             64267 when "00001100001010",
                             64185 when "00001100001011",
                             64103 when "00001100001100",
                             64020 when "00001100001101",
                             63939 when "00001100001110",
                             63857 when "00001100001111",
                             63776 when "00001100010000",
                             63694 when "00001100010001",
                             63613 when "00001100010010",
                             63532 when "00001100010011",
                             63452 when "00001100010100",
                             63371 when "00001100010101",
                             63291 when "00001100010110",
                             63211 when "00001100010111",
                             63131 when "00001100011000",
                             63052 when "00001100011001",
                             62972 when "00001100011010",
                             62893 when "00001100011011",
                             62814 when "00001100011100",
                             62735 when "00001100011101",
                             62657 when "00001100011110",
                             62578 when "00001100011111",
                             62500 when "00001100100000",
                             62422 when "00001100100001",
                             62344 when "00001100100010",
                             62267 when "00001100100011",
                             62189 when "00001100100100",
                             62112 when "00001100100101",
                             62035 when "00001100100110",
                             61958 when "00001100100111",
                             61881 when "00001100101000",
                             61805 when "00001100101001",
                             61728 when "00001100101010",
                             61652 when "00001100101011",
                             61576 when "00001100101100",
                             61501 when "00001100101101",
                             61425 when "00001100101110",
                             61350 when "00001100101111",
                             61275 when "00001100110000",
                             61200 when "00001100110001",
                             61125 when "00001100110010",
                             61050 when "00001100110011",
                             60976 when "00001100110100",
                             60901 when "00001100110101",
                             60827 when "00001100110110",
                             60753 when "00001100110111",
                             60680 when "00001100111000",
                             60606 when "00001100111001",
                             60533 when "00001100111010",
                             60459 when "00001100111011",
                             60386 when "00001100111100",
                             60314 when "00001100111101",
                             60241 when "00001100111110",
                             60168 when "00001100111111",
                             60096 when "00001101000000",
                             60024 when "00001101000001",
                             59952 when "00001101000010",
                             59880 when "00001101000011",
                             59809 when "00001101000100",
                             59737 when "00001101000101",
                             59666 when "00001101000110",
                             59595 when "00001101000111",
                             59524 when "00001101001000",
                             59453 when "00001101001001",
                             59382 when "00001101001010",
                             59312 when "00001101001011",
                             59242 when "00001101001100",
                             59172 when "00001101001101",
                             59102 when "00001101001110",
                             59032 when "00001101001111",
                             58962 when "00001101010000",
                             58893 when "00001101010001",
                             58824 when "00001101010010",
                             58754 when "00001101010011",
                             58685 when "00001101010100",
                             58617 when "00001101010101",
                             58548 when "00001101010110",
                             58480 when "00001101010111",
                             58411 when "00001101011000",
                             58343 when "00001101011001",
                             58275 when "00001101011010",
                             58207 when "00001101011011",
                             58140 when "00001101011100",
                             58072 when "00001101011101",
                             58005 when "00001101011110",
                             57937 when "00001101011111",
                             57870 when "00001101100000",
                             57803 when "00001101100001",
                             57737 when "00001101100010",
                             57670 when "00001101100011",
                             57604 when "00001101100100",
                             57537 when "00001101100101",
                             57471 when "00001101100110",
                             57405 when "00001101100111",
                             57339 when "00001101101000",
                             57274 when "00001101101001",
                             57208 when "00001101101010",
                             57143 when "00001101101011",
                             57078 when "00001101101100",
                             57013 when "00001101101101",
                             56948 when "00001101101110",
                             56883 when "00001101101111",
                             56818 when "00001101110000",
                             56754 when "00001101110001",
                             56689 when "00001101110010",
                             56625 when "00001101110011",
                             56561 when "00001101110100",
                             56497 when "00001101110101",
                             56433 when "00001101110110",
                             56370 when "00001101110111",
                             56306 when "00001101111000",
                             56243 when "00001101111001",
                             56180 when "00001101111010",
                             56117 when "00001101111011",
                             56054 when "00001101111100",
                             55991 when "00001101111101",
                             55928 when "00001101111110",
                             55866 when "00001101111111",
                             55804 when "00001110000000",
                             55741 when "00001110000001",
                             55679 when "00001110000010",
                             55617 when "00001110000011",
                             55556 when "00001110000100",
                             55494 when "00001110000101",
                             55432 when "00001110000110",
                             55371 when "00001110000111",
                             55310 when "00001110001000",
                             55249 when "00001110001001",
                             55188 when "00001110001010",
                             55127 when "00001110001011",
                             55066 when "00001110001100",
                             55006 when "00001110001101",
                             54945 when "00001110001110",
                             54885 when "00001110001111",
                             54825 when "00001110010000",
                             54765 when "00001110010001",
                             54705 when "00001110010010",
                             54645 when "00001110010011",
                             54585 when "00001110010100",
                             54526 when "00001110010101",
                             54466 when "00001110010110",
                             54407 when "00001110010111",
                             54348 when "00001110011000",
                             54289 when "00001110011001",
                             54230 when "00001110011010",
                             54171 when "00001110011011",
                             54113 when "00001110011100",
                             54054 when "00001110011101",
                             53996 when "00001110011110",
                             53937 when "00001110011111",
                             53879 when "00001110100000",
                             53821 when "00001110100001",
                             53763 when "00001110100010",
                             53706 when "00001110100011",
                             53648 when "00001110100100",
                             53591 when "00001110100101",
                             53533 when "00001110100110",
                             53476 when "00001110100111",
                             53419 when "00001110101000",
                             53362 when "00001110101001",
                             53305 when "00001110101010",
                             53248 when "00001110101011",
                             53191 when "00001110101100",
                             53135 when "00001110101101",
                             53079 when "00001110101110",
                             53022 when "00001110101111",
                             52966 when "00001110110000",
                             52910 when "00001110110001",
                             52854 when "00001110110010",
                             52798 when "00001110110011",
                             52743 when "00001110110100",
                             52687 when "00001110110101",
                             52632 when "00001110110110",
                             52576 when "00001110110111",
                             52521 when "00001110111000",
                             52466 when "00001110111001",
                             52411 when "00001110111010",
                             52356 when "00001110111011",
                             52301 when "00001110111100",
                             52247 when "00001110111101",
                             52192 when "00001110111110",
                             52138 when "00001110111111",
                             52083 when "00001111000000",
                             52029 when "00001111000001",
                             51975 when "00001111000010",
                             51921 when "00001111000011",
                             51867 when "00001111000100",
                             51813 when "00001111000101",
                             51760 when "00001111000110",
                             51706 when "00001111000111",
                             51653 when "00001111001000",
                             51600 when "00001111001001",
                             51546 when "00001111001010",
                             51493 when "00001111001011",
                             51440 when "00001111001100",
                             51387 when "00001111001101",
                             51335 when "00001111001110",
                             51282 when "00001111001111",
                             51230 when "00001111010000",
                             51177 when "00001111010001",
                             51125 when "00001111010010",
                             51073 when "00001111010011",
                             51020 when "00001111010100",
                             50968 when "00001111010101",
                             50916 when "00001111010110",
                             50865 when "00001111010111",
                             50813 when "00001111011000",
                             50761 when "00001111011001",
                             50710 when "00001111011010",
                             50659 when "00001111011011",
                             50607 when "00001111011100",
                             50556 when "00001111011101",
                             50505 when "00001111011110",
                             50454 when "00001111011111",
                             50403 when "00001111100000",
                             50352 when "00001111100001",
                             50302 when "00001111100010",
                             50251 when "00001111100011",
                             50201 when "00001111100100",
                             50150 when "00001111100101",
                             50100 when "00001111100110",
                             50050 when "00001111100111",
                             50000 when "00001111101000",
                             49950 when "00001111101001",
                             49900 when "00001111101010",
                             49850 when "00001111101011",
                             49801 when "00001111101100",
                             49751 when "00001111101101",
                             49702 when "00001111101110",
                             49652 when "00001111101111",
                             49603 when "00001111110000",
                             49554 when "00001111110001",
                             49505 when "00001111110010",
                             49456 when "00001111110011",
                             49407 when "00001111110100",
                             49358 when "00001111110101",
                             49310 when "00001111110110",
                             49261 when "00001111110111",
                             49213 when "00001111111000",
                             49164 when "00001111111001",
                             49116 when "00001111111010",
                             49068 when "00001111111011",
                             49020 when "00001111111100",
                             48972 when "00001111111101",
                             48924 when "00001111111110",
                             48876 when "00001111111111",
                             48828 when "00010000000000",
                             48780 when "00010000000001",
                             48733 when "00010000000010",
                             48685 when "00010000000011",
                             48638 when "00010000000100",
                             48591 when "00010000000101",
                             48544 when "00010000000110",
                             48497 when "00010000000111",
                             48450 when "00010000001000",
                             48403 when "00010000001001",
                             48356 when "00010000001010",
                             48309 when "00010000001011",
                             48263 when "00010000001100",
                             48216 when "00010000001101",
                             48170 when "00010000001110",
                             48123 when "00010000001111",
                             48077 when "00010000010000",
                             48031 when "00010000010001",
                             47985 when "00010000010010",
                             47939 when "00010000010011",
                             47893 when "00010000010100",
                             47847 when "00010000010101",
                             47801 when "00010000010110",
                             47755 when "00010000010111",
                             47710 when "00010000011000",
                             47664 when "00010000011001",
                             47619 when "00010000011010",
                             47574 when "00010000011011",
                             47529 when "00010000011100",
                             47483 when "00010000011101",
                             47438 when "00010000011110",
                             47393 when "00010000011111",
                             47348 when "00010000100000",
                             47304 when "00010000100001",
                             47259 when "00010000100010",
                             47214 when "00010000100011",
                             47170 when "00010000100100",
                             47125 when "00010000100101",
                             47081 when "00010000100110",
                             47037 when "00010000100111",
                             46992 when "00010000101000",
                             46948 when "00010000101001",
                             46904 when "00010000101010",
                             46860 when "00010000101011",
                             46816 when "00010000101100",
                             46773 when "00010000101101",
                             46729 when "00010000101110",
                             46685 when "00010000101111",
                             46642 when "00010000110000",
                             46598 when "00010000110001",
                             46555 when "00010000110010",
                             46512 when "00010000110011",
                             46468 when "00010000110100",
                             46425 when "00010000110101",
                             46382 when "00010000110110",
                             46339 when "00010000110111",
                             46296 when "00010000111000",
                             46253 when "00010000111001",
                             46211 when "00010000111010",
                             46168 when "00010000111011",
                             46125 when "00010000111100",
                             46083 when "00010000111101",
                             46041 when "00010000111110",
                             45998 when "00010000111111",
                             45956 when "00010001000000",
                             45914 when "00010001000001",
                             45872 when "00010001000010",
                             45830 when "00010001000011",
                             45788 when "00010001000100",
                             45746 when "00010001000101",
                             45704 when "00010001000110",
                             45662 when "00010001000111",
                             45620 when "00010001001000",
                             45579 when "00010001001001",
                             45537 when "00010001001010",
                             45496 when "00010001001011",
                             45455 when "00010001001100",
                             45413 when "00010001001101",
                             45372 when "00010001001110",
                             45331 when "00010001001111",
                             45290 when "00010001010000",
                             45249 when "00010001010001",
                             45208 when "00010001010010",
                             45167 when "00010001010011",
                             45126 when "00010001010100",
                             45086 when "00010001010101",
                             45045 when "00010001010110",
                             45005 when "00010001010111",
                             44964 when "00010001011000",
                             44924 when "00010001011001",
                             44883 when "00010001011010",
                             44843 when "00010001011011",
                             44803 when "00010001011100",
                             44763 when "00010001011101",
                             44723 when "00010001011110",
                             44683 when "00010001011111",
                             44643 when "00010001100000",
                             44603 when "00010001100001",
                             44563 when "00010001100010",
                             44524 when "00010001100011",
                             44484 when "00010001100100",
                             44444 when "00010001100101",
                             44405 when "00010001100110",
                             44366 when "00010001100111",
                             44326 when "00010001101000",
                             44287 when "00010001101001",
                             44248 when "00010001101010",
                             44209 when "00010001101011",
                             44170 when "00010001101100",
                             44131 when "00010001101101",
                             44092 when "00010001101110",
                             44053 when "00010001101111",
                             44014 when "00010001110000",
                             43975 when "00010001110001",
                             43937 when "00010001110010",
                             43898 when "00010001110011",
                             43860 when "00010001110100",
                             43821 when "00010001110101",
                             43783 when "00010001110110",
                             43745 when "00010001110111",
                             43706 when "00010001111000",
                             43668 when "00010001111001",
                             43630 when "00010001111010",
                             43592 when "00010001111011",
                             43554 when "00010001111100",
                             43516 when "00010001111101",
                             43478 when "00010001111110",
                             43440 when "00010001111111",
                             43403 when "00010010000000",
                             43365 when "00010010000001",
                             43328 when "00010010000010",
                             43290 when "00010010000011",
                             43253 when "00010010000100",
                             43215 when "00010010000101",
                             43178 when "00010010000110",
                             43141 when "00010010000111",
                             43103 when "00010010001000",
                             43066 when "00010010001001",
                             43029 when "00010010001010",
                             42992 when "00010010001011",
                             42955 when "00010010001100",
                             42918 when "00010010001101",
                             42882 when "00010010001110",
                             42845 when "00010010001111",
                             42808 when "00010010010000",
                             42772 when "00010010010001",
                             42735 when "00010010010010",
                             42699 when "00010010010011",
                             42662 when "00010010010100",
                             42626 when "00010010010101",
                             42589 when "00010010010110",
                             42553 when "00010010010111",
                             42517 when "00010010011000",
                             42481 when "00010010011001",
                             42445 when "00010010011010",
                             42409 when "00010010011011",
                             42373 when "00010010011100",
                             42337 when "00010010011101",
                             42301 when "00010010011110",
                             42265 when "00010010011111",
                             42230 when "00010010100000",
                             42194 when "00010010100001",
                             42159 when "00010010100010",
                             42123 when "00010010100011",
                             42088 when "00010010100100",
                             42052 when "00010010100101",
                             42017 when "00010010100110",
                             41982 when "00010010100111",
                             41946 when "00010010101000",
                             41911 when "00010010101001",
                             41876 when "00010010101010",
                             41841 when "00010010101011",
                             41806 when "00010010101100",
                             41771 when "00010010101101",
                             41736 when "00010010101110",
                             41701 when "00010010101111",
                             41667 when "00010010110000",
                             41632 when "00010010110001",
                             41597 when "00010010110010",
                             41563 when "00010010110011",
                             41528 when "00010010110100",
                             41494 when "00010010110101",
                             41459 when "00010010110110",
                             41425 when "00010010110111",
                             41391 when "00010010111000",
                             41356 when "00010010111001",
                             41322 when "00010010111010",
                             41288 when "00010010111011",
                             41254 when "00010010111100",
                             41220 when "00010010111101",
                             41186 when "00010010111110",
                             41152 when "00010010111111",
                             41118 when "00010011000000",
                             41085 when "00010011000001",
                             41051 when "00010011000010",
                             41017 when "00010011000011",
                             40984 when "00010011000100",
                             40950 when "00010011000101",
                             40917 when "00010011000110",
                             40883 when "00010011000111",
                             40850 when "00010011001000",
                             40816 when "00010011001001",
                             40783 when "00010011001010",
                             40750 when "00010011001011",
                             40717 when "00010011001100",
                             40683 when "00010011001101",
                             40650 when "00010011001110",
                             40617 when "00010011001111",
                             40584 when "00010011010000",
                             40552 when "00010011010001",
                             40519 when "00010011010010",
                             40486 when "00010011010011",
                             40453 when "00010011010100",
                             40420 when "00010011010101",
                             40388 when "00010011010110",
                             40355 when "00010011010111",
                             40323 when "00010011011000",
                             40290 when "00010011011001",
                             40258 when "00010011011010",
                             40225 when "00010011011011",
                             40193 when "00010011011100",
                             40161 when "00010011011101",
                             40128 when "00010011011110",
                             40096 when "00010011011111",
                             40064 when "00010011100000",
                             40032 when "00010011100001",
                             40000 when "00010011100010",
                             39968 when "00010011100011",
                             39936 when "00010011100100",
                             39904 when "00010011100101",
                             39872 when "00010011100110",
                             39841 when "00010011100111",
                             39809 when "00010011101000",
                             39777 when "00010011101001",
                             39746 when "00010011101010",
                             39714 when "00010011101011",
                             39683 when "00010011101100",
                             39651 when "00010011101101",
                             39620 when "00010011101110",
                             39588 when "00010011101111",
                             39557 when "00010011110000",
                             39526 when "00010011110001",
                             39494 when "00010011110010",
                             39463 when "00010011110011",
                             39432 when "00010011110100",
                             39401 when "00010011110101",
                             39370 when "00010011110110",
                             39339 when "00010011110111",
                             39308 when "00010011111000",
                             39277 when "00010011111001",
                             39246 when "00010011111010",
                             39216 when "00010011111011",
                             39185 when "00010011111100",
                             39154 when "00010011111101",
                             39124 when "00010011111110",
                             39093 when "00010011111111",
                             39063 when "00010100000000",
                             39032 when "00010100000001",
                             39002 when "00010100000010",
                             38971 when "00010100000011",
                             38941 when "00010100000100",
                             38911 when "00010100000101",
                             38880 when "00010100000110",
                             38850 when "00010100000111",
                             38820 when "00010100001000",
                             38790 when "00010100001001",
                             38760 when "00010100001010",
                             38730 when "00010100001011",
                             38700 when "00010100001100",
                             38670 when "00010100001101",
                             38640 when "00010100001110",
                             38610 when "00010100001111",
                             38580 when "00010100010000",
                             38551 when "00010100010001",
                             38521 when "00010100010010",
                             38491 when "00010100010011",
                             38462 when "00010100010100",
                             38432 when "00010100010101",
                             38402 when "00010100010110",
                             38373 when "00010100010111",
                             38344 when "00010100011000",
                             38314 when "00010100011001",
                             38285 when "00010100011010",
                             38256 when "00010100011011",
                             38226 when "00010100011100",
                             38197 when "00010100011101",
                             38168 when "00010100011110",
                             38139 when "00010100011111",
                             38110 when "00010100100000",
                             38081 when "00010100100001",
                             38052 when "00010100100010",
                             38023 when "00010100100011",
                             37994 when "00010100100100",
                             37965 when "00010100100101",
                             37936 when "00010100100110",
                             37908 when "00010100100111",
                             37879 when "00010100101000",
                             37850 when "00010100101001",
                             37821 when "00010100101010",
                             37793 when "00010100101011",
                             37764 when "00010100101100",
                             37736 when "00010100101101",
                             37707 when "00010100101110",
                             37679 when "00010100101111",
                             37651 when "00010100110000",
                             37622 when "00010100110001",
                             37594 when "00010100110010",
                             37566 when "00010100110011",
                             37538 when "00010100110100",
                             37509 when "00010100110101",
                             37481 when "00010100110110",
                             37453 when "00010100110111",
                             37425 when "00010100111000",
                             37397 when "00010100111001",
                             37369 when "00010100111010",
                             37341 when "00010100111011",
                             37313 when "00010100111100",
                             37286 when "00010100111101",
                             37258 when "00010100111110",
                             37230 when "00010100111111",
                             37202 when "00010101000000",
                             37175 when "00010101000001",
                             37147 when "00010101000010",
                             37120 when "00010101000011",
                             37092 when "00010101000100",
                             37064 when "00010101000101",
                             37037 when "00010101000110",
                             37010 when "00010101000111",
                             36982 when "00010101001000",
                             36955 when "00010101001001",
                             36928 when "00010101001010",
                             36900 when "00010101001011",
                             36873 when "00010101001100",
                             36846 when "00010101001101",
                             36819 when "00010101001110",
                             36792 when "00010101001111",
                             36765 when "00010101010000",
                             36738 when "00010101010001",
                             36711 when "00010101010010",
                             36684 when "00010101010011",
                             36657 when "00010101010100",
                             36630 when "00010101010101",
                             36603 when "00010101010110",
                             36576 when "00010101010111",
                             36550 when "00010101011000",
                             36523 when "00010101011001",
                             36496 when "00010101011010",
                             36470 when "00010101011011",
                             36443 when "00010101011100",
                             36417 when "00010101011101",
                             36390 when "00010101011110",
                             36364 when "00010101011111",
                             36337 when "00010101100000",
                             36311 when "00010101100001",
                             36284 when "00010101100010",
                             36258 when "00010101100011",
                             36232 when "00010101100100",
                             36206 when "00010101100101",
                             36179 when "00010101100110",
                             36153 when "00010101100111",
                             36127 when "00010101101000",
                             36101 when "00010101101001",
                             36075 when "00010101101010",
                             36049 when "00010101101011",
                             36023 when "00010101101100",
                             35997 when "00010101101101",
                             35971 when "00010101101110",
                             35945 when "00010101101111",
                             35920 when "00010101110000",
                             35894 when "00010101110001",
                             35868 when "00010101110010",
                             35842 when "00010101110011",
                             35817 when "00010101110100",
                             35791 when "00010101110101",
                             35765 when "00010101110110",
                             35740 when "00010101110111",
                             35714 when "00010101111000",
                             35689 when "00010101111001",
                             35663 when "00010101111010",
                             35638 when "00010101111011",
                             35613 when "00010101111100",
                             35587 when "00010101111101",
                             35562 when "00010101111110",
                             35537 when "00010101111111",
                             35511 when "00010110000000",
                             35486 when "00010110000001",
                             35461 when "00010110000010",
                             35436 when "00010110000011",
                             35411 when "00010110000100",
                             35386 when "00010110000101",
                             35361 when "00010110000110",
                             35336 when "00010110000111",
                             35311 when "00010110001000",
                             35286 when "00010110001001",
                             35261 when "00010110001010",
                             35236 when "00010110001011",
                             35211 when "00010110001100",
                             35186 when "00010110001101",
                             35162 when "00010110001110",
                             35137 when "00010110001111",
                             35112 when "00010110010000",
                             35088 when "00010110010001",
                             35063 when "00010110010010",
                             35039 when "00010110010011",
                             35014 when "00010110010100",
                             34990 when "00010110010101",
                             34965 when "00010110010110",
                             34941 when "00010110010111",
                             34916 when "00010110011000",
                             34892 when "00010110011001",
                             34868 when "00010110011010",
                             34843 when "00010110011011",
                             34819 when "00010110011100",
                             34795 when "00010110011101",
                             34771 when "00010110011110",
                             34746 when "00010110011111",
                             34722 when "00010110100000",
                             34698 when "00010110100001",
                             34674 when "00010110100010",
                             34650 when "00010110100011",
                             34626 when "00010110100100",
                             34602 when "00010110100101",
                             34578 when "00010110100110",
                             34554 when "00010110100111",
                             34530 when "00010110101000",
                             34507 when "00010110101001",
                             34483 when "00010110101010",
                             34459 when "00010110101011",
                             34435 when "00010110101100",
                             34412 when "00010110101101",
                             34388 when "00010110101110",
                             34364 when "00010110101111",
                             34341 when "00010110110000",
                             34317 when "00010110110001",
                             34294 when "00010110110010",
                             34270 when "00010110110011",
                             34247 when "00010110110100",
                             34223 when "00010110110101",
                             34200 when "00010110110110",
                             34176 when "00010110110111",
                             34153 when "00010110111000",
                             34130 when "00010110111001",
                             34106 when "00010110111010",
                             34083 when "00010110111011",
                             34060 when "00010110111100",
                             34037 when "00010110111101",
                             34014 when "00010110111110",
                             33990 when "00010110111111",
                             33967 when "00010111000000",
                             33944 when "00010111000001",
                             33921 when "00010111000010",
                             33898 when "00010111000011",
                             33875 when "00010111000100",
                             33852 when "00010111000101",
                             33829 when "00010111000110",
                             33807 when "00010111000111",
                             33784 when "00010111001000",
                             33761 when "00010111001001",
                             33738 when "00010111001010",
                             33715 when "00010111001011",
                             33693 when "00010111001100",
                             33670 when "00010111001101",
                             33647 when "00010111001110",
                             33625 when "00010111001111",
                             33602 when "00010111010000",
                             33580 when "00010111010001",
                             33557 when "00010111010010",
                             33535 when "00010111010011",
                             33512 when "00010111010100",
                             33490 when "00010111010101",
                             33467 when "00010111010110",
                             33445 when "00010111010111",
                             33422 when "00010111011000",
                             33400 when "00010111011001",
                             33378 when "00010111011010",
                             33356 when "00010111011011",
                             33333 when "00010111011100",
                             33311 when "00010111011101",
                             33289 when "00010111011110",
                             33267 when "00010111011111",
                             33245 when "00010111100000",
                             33223 when "00010111100001",
                             33201 when "00010111100010",
                             33179 when "00010111100011",
                             33156 when "00010111100100",
                             33135 when "00010111100101",
                             33113 when "00010111100110",
                             33091 when "00010111100111",
                             33069 when "00010111101000",
                             33047 when "00010111101001",
                             33025 when "00010111101010",
                             33003 when "00010111101011",
                             32982 when "00010111101100",
                             32960 when "00010111101101",
                             32938 when "00010111101110",
                             32916 when "00010111101111",
                             32895 when "00010111110000",
                             32873 when "00010111110001",
                             32852 when "00010111110010",
                             32830 when "00010111110011",
                             32808 when "00010111110100",
                             32787 when "00010111110101",
                             32765 when "00010111110110",
                             32744 when "00010111110111",
                             32723 when "00010111111000",
                             32701 when "00010111111001",
                             32680 when "00010111111010",
                             32658 when "00010111111011",
                             32637 when "00010111111100",
                             32616 when "00010111111101",
                             32595 when "00010111111110",
                             32573 when "00010111111111",
                             32552 when "00011000000000",
                             32531 when "00011000000001",
                             32510 when "00011000000010",
                             32489 when "00011000000011",
                             32468 when "00011000000100",
                             32446 when "00011000000101",
                             32425 when "00011000000110",
                             32404 when "00011000000111",
                             32383 when "00011000001000",
                             32362 when "00011000001001",
                             32342 when "00011000001010",
                             32321 when "00011000001011",
                             32300 when "00011000001100",
                             32279 when "00011000001101",
                             32258 when "00011000001110",
                             32237 when "00011000001111",
                             32216 when "00011000010000",
                             32196 when "00011000010001",
                             32175 when "00011000010010",
                             32154 when "00011000010011",
                             32134 when "00011000010100",
                             32113 when "00011000010101",
                             32092 when "00011000010110",
                             32072 when "00011000010111",
                             32051 when "00011000011000",
                             32031 when "00011000011001",
                             32010 when "00011000011010",
                             31990 when "00011000011011",
                             31969 when "00011000011100",
                             31949 when "00011000011101",
                             31928 when "00011000011110",
                             31908 when "00011000011111",
                             31888 when "00011000100000",
                             31867 when "00011000100001",
                             31847 when "00011000100010",
                             31827 when "00011000100011",
                             31807 when "00011000100100",
                             31786 when "00011000100101",
                             31766 when "00011000100110",
                             31746 when "00011000100111",
                             31726 when "00011000101000",
                             31706 when "00011000101001",
                             31686 when "00011000101010",
                             31666 when "00011000101011",
                             31646 when "00011000101100",
                             31626 when "00011000101101",
                             31606 when "00011000101110",
                             31586 when "00011000101111",
                             31566 when "00011000110000",
                             31546 when "00011000110001",
                             31526 when "00011000110010",
                             31506 when "00011000110011",
                             31486 when "00011000110100",
                             31466 when "00011000110101",
                             31447 when "00011000110110",
                             31427 when "00011000110111",
                             31407 when "00011000111000",
                             31387 when "00011000111001",
                             31368 when "00011000111010",
                             31348 when "00011000111011",
                             31328 when "00011000111100",
                             31309 when "00011000111101",
                             31289 when "00011000111110",
                             31270 when "00011000111111",
                             31250 when "00011001000000",
                             31230 when "00011001000001",
                             31211 when "00011001000010",
                             31192 when "00011001000011",
                             31172 when "00011001000100",
                             31153 when "00011001000101",
                             31133 when "00011001000110",
                             31114 when "00011001000111",
                             31095 when "00011001001000",
                             31075 when "00011001001001",
                             31056 when "00011001001010",
                             31037 when "00011001001011",
                             31017 when "00011001001100",
                             30998 when "00011001001101",
                             30979 when "00011001001110",
                             30960 when "00011001001111",
                             30941 when "00011001010000",
                             30921 when "00011001010001",
                             30902 when "00011001010010",
                             30883 when "00011001010011",
                             30864 when "00011001010100",
                             30845 when "00011001010101",
                             30826 when "00011001010110",
                             30807 when "00011001010111",
                             30788 when "00011001011000",
                             30769 when "00011001011001",
                             30750 when "00011001011010",
                             30731 when "00011001011011",
                             30713 when "00011001011100",
                             30694 when "00011001011101",
                             30675 when "00011001011110",
                             30656 when "00011001011111",
                             30637 when "00011001100000",
                             30618 when "00011001100001",
                             30600 when "00011001100010",
                             30581 when "00011001100011",
                             30562 when "00011001100100",
                             30544 when "00011001100101",
                             30525 when "00011001100110",
                             30506 when "00011001100111",
                             30488 when "00011001101000",
                             30469 when "00011001101001",
                             30451 when "00011001101010",
                             30432 when "00011001101011",
                             30414 when "00011001101100",
                             30395 when "00011001101101",
                             30377 when "00011001101110",
                             30358 when "00011001101111",
                             30340 when "00011001110000",
                             30321 when "00011001110001",
                             30303 when "00011001110010",
                             30285 when "00011001110011",
                             30266 when "00011001110100",
                             30248 when "00011001110101",
                             30230 when "00011001110110",
                             30211 when "00011001110111",
                             30193 when "00011001111000",
                             30175 when "00011001111001",
                             30157 when "00011001111010",
                             30139 when "00011001111011",
                             30120 when "00011001111100",
                             30102 when "00011001111101",
                             30084 when "00011001111110",
                             30066 when "00011001111111",
                             30048 when "00011010000000",
                             30030 when "00011010000001",
                             30012 when "00011010000010",
                             29994 when "00011010000011",
                             29976 when "00011010000100",
                             29958 when "00011010000101",
                             29940 when "00011010000110",
                             29922 when "00011010000111",
                             29904 when "00011010001000",
                             29886 when "00011010001001",
                             29869 when "00011010001010",
                             29851 when "00011010001011",
                             29833 when "00011010001100",
                             29815 when "00011010001101",
                             29797 when "00011010001110",
                             29780 when "00011010001111",
                             29762 when "00011010010000",
                             29744 when "00011010010001",
                             29727 when "00011010010010",
                             29709 when "00011010010011",
                             29691 when "00011010010100",
                             29674 when "00011010010101",
                             29656 when "00011010010110",
                             29638 when "00011010010111",
                             29621 when "00011010011000",
                             29603 when "00011010011001",
                             29586 when "00011010011010",
                             29568 when "00011010011011",
                             29551 when "00011010011100",
                             29533 when "00011010011101",
                             29516 when "00011010011110",
                             29499 when "00011010011111",
                             29481 when "00011010100000",
                             29464 when "00011010100001",
                             29446 when "00011010100010",
                             29429 when "00011010100011",
                             29412 when "00011010100100",
                             29394 when "00011010100101",
                             29377 when "00011010100110",
                             29360 when "00011010100111",
                             29343 when "00011010101000",
                             29326 when "00011010101001",
                             29308 when "00011010101010",
                             29291 when "00011010101011",
                             29274 when "00011010101100",
                             29257 when "00011010101101",
                             29240 when "00011010101110",
                             29223 when "00011010101111",
                             29206 when "00011010110000",
                             29189 when "00011010110001",
                             29172 when "00011010110010",
                             29155 when "00011010110011",
                             29138 when "00011010110100",
                             29121 when "00011010110101",
                             29104 when "00011010110110",
                             29087 when "00011010110111",
                             29070 when "00011010111000",
                             29053 when "00011010111001",
                             29036 when "00011010111010",
                             29019 when "00011010111011",
                             29002 when "00011010111100",
                             28986 when "00011010111101",
                             28969 when "00011010111110",
                             28952 when "00011010111111",
                             28935 when "00011011000000",
                             28918 when "00011011000001",
                             28902 when "00011011000010",
                             28885 when "00011011000011",
                             28868 when "00011011000100",
                             28852 when "00011011000101",
                             28835 when "00011011000110",
                             28818 when "00011011000111",
                             28802 when "00011011001000",
                             28785 when "00011011001001",
                             28769 when "00011011001010",
                             28752 when "00011011001011",
                             28736 when "00011011001100",
                             28719 when "00011011001101",
                             28703 when "00011011001110",
                             28686 when "00011011001111",
                             28670 when "00011011010000",
                             28653 when "00011011010001",
                             28637 when "00011011010010",
                             28620 when "00011011010011",
                             28604 when "00011011010100",
                             28588 when "00011011010101",
                             28571 when "00011011010110",
                             28555 when "00011011010111",
                             28539 when "00011011011000",
                             28523 when "00011011011001",
                             28506 when "00011011011010",
                             28490 when "00011011011011",
                             28474 when "00011011011100",
                             28458 when "00011011011101",
                             28441 when "00011011011110",
                             28425 when "00011011011111",
                             28409 when "00011011100000",
                             28393 when "00011011100001",
                             28377 when "00011011100010",
                             28361 when "00011011100011",
                             28345 when "00011011100100",
                             28329 when "00011011100101",
                             28313 when "00011011100110",
                             28297 when "00011011100111",
                             28281 when "00011011101000",
                             28265 when "00011011101001",
                             28249 when "00011011101010",
                             28233 when "00011011101011",
                             28217 when "00011011101100",
                             28201 when "00011011101101",
                             28185 when "00011011101110",
                             28169 when "00011011101111",
                             28153 when "00011011110000",
                             28137 when "00011011110001",
                             28121 when "00011011110010",
                             28106 when "00011011110011",
                             28090 when "00011011110100",
                             28074 when "00011011110101",
                             28058 when "00011011110110",
                             28043 when "00011011110111",
                             28027 when "00011011111000",
                             28011 when "00011011111001",
                             27996 when "00011011111010",
                             27980 when "00011011111011",
                             27964 when "00011011111100",
                             27949 when "00011011111101",
                             27933 when "00011011111110",
                             27917 when "00011011111111",
                             27902 when "00011100000000",
                             27886 when "00011100000001",
                             27871 when "00011100000010",
                             27855 when "00011100000011",
                             27840 when "00011100000100",
                             27824 when "00011100000101",
                             27809 when "00011100000110",
                             27793 when "00011100000111",
                             27778 when "00011100001000",
                             27762 when "00011100001001",
                             27747 when "00011100001010",
                             27732 when "00011100001011",
                             27716 when "00011100001100",
                             27701 when "00011100001101",
                             27685 when "00011100001110",
                             27670 when "00011100001111",
                             27655 when "00011100010000",
                             27640 when "00011100010001",
                             27624 when "00011100010010",
                             27609 when "00011100010011",
                             27594 when "00011100010100",
                             27579 when "00011100010101",
                             27563 when "00011100010110",
                             27548 when "00011100010111",
                             27533 when "00011100011000",
                             27518 when "00011100011001",
                             27503 when "00011100011010",
                             27488 when "00011100011011",
                             27473 when "00011100011100",
                             27457 when "00011100011101",
                             27442 when "00011100011110",
                             27427 when "00011100011111",
                             27412 when "00011100100000",
                             27397 when "00011100100001",
                             27382 when "00011100100010",
                             27367 when "00011100100011",
                             27352 when "00011100100100",
                             27337 when "00011100100101",
                             27322 when "00011100100110",
                             27307 when "00011100100111",
                             27293 when "00011100101000",
                             27278 when "00011100101001",
                             27263 when "00011100101010",
                             27248 when "00011100101011",
                             27233 when "00011100101100",
                             27218 when "00011100101101",
                             27203 when "00011100101110",
                             27189 when "00011100101111",
                             27174 when "00011100110000",
                             27159 when "00011100110001",
                             27144 when "00011100110010",
                             27130 when "00011100110011",
                             27115 when "00011100110100",
                             27100 when "00011100110101",
                             27086 when "00011100110110",
                             27071 when "00011100110111",
                             27056 when "00011100111000",
                             27042 when "00011100111001",
                             27027 when "00011100111010",
                             27012 when "00011100111011",
                             26998 when "00011100111100",
                             26983 when "00011100111101",
                             26969 when "00011100111110",
                             26954 when "00011100111111",
                             26940 when "00011101000000",
                             26925 when "00011101000001",
                             26911 when "00011101000010",
                             26896 when "00011101000011",
                             26882 when "00011101000100",
                             26867 when "00011101000101",
                             26853 when "00011101000110",
                             26838 when "00011101000111",
                             26824 when "00011101001000",
                             26810 when "00011101001001",
                             26795 when "00011101001010",
                             26781 when "00011101001011",
                             26767 when "00011101001100",
                             26752 when "00011101001101",
                             26738 when "00011101001110",
                             26724 when "00011101001111",
                             26709 when "00011101010000",
                             26695 when "00011101010001",
                             26681 when "00011101010010",
                             26667 when "00011101010011",
                             26652 when "00011101010100",
                             26638 when "00011101010101",
                             26624 when "00011101010110",
                             26610 when "00011101010111",
                             26596 when "00011101011000",
                             26582 when "00011101011001",
                             26567 when "00011101011010",
                             26553 when "00011101011011",
                             26539 when "00011101011100",
                             26525 when "00011101011101",
                             26511 when "00011101011110",
                             26497 when "00011101011111",
                             26483 when "00011101100000",
                             26469 when "00011101100001",
                             26455 when "00011101100010",
                             26441 when "00011101100011",
                             26427 when "00011101100100",
                             26413 when "00011101100101",
                             26399 when "00011101100110",
                             26385 when "00011101100111",
                             26371 when "00011101101000",
                             26357 when "00011101101001",
                             26344 when "00011101101010",
                             26330 when "00011101101011",
                             26316 when "00011101101100",
                             26302 when "00011101101101",
                             26288 when "00011101101110",
                             26274 when "00011101101111",
                             26261 when "00011101110000",
                             26247 when "00011101110001",
                             26233 when "00011101110010",
                             26219 when "00011101110011",
                             26205 when "00011101110100",
                             26192 when "00011101110101",
                             26178 when "00011101110110",
                             26164 when "00011101110111",
                             26151 when "00011101111000",
                             26137 when "00011101111001",
                             26123 when "00011101111010",
                             26110 when "00011101111011",
                             26096 when "00011101111100",
                             26082 when "00011101111101",
                             26069 when "00011101111110",
                             26055 when "00011101111111",
                             26042 when "00011110000000",
                             26028 when "00011110000001",
                             26015 when "00011110000010",
                             26001 when "00011110000011",
                             25988 when "00011110000100",
                             25974 when "00011110000101",
                             25961 when "00011110000110",
                             25947 when "00011110000111",
                             25934 when "00011110001000",
                             25920 when "00011110001001",
                             25907 when "00011110001010",
                             25893 when "00011110001011",
                             25880 when "00011110001100",
                             25867 when "00011110001101",
                             25853 when "00011110001110",
                             25840 when "00011110001111",
                             25826 when "00011110010000",
                             25813 when "00011110010001",
                             25800 when "00011110010010",
                             25786 when "00011110010011",
                             25773 when "00011110010100",
                             25760 when "00011110010101",
                             25747 when "00011110010110",
                             25733 when "00011110010111",
                             25720 when "00011110011000",
                             25707 when "00011110011001",
                             25694 when "00011110011010",
                             25681 when "00011110011011",
                             25667 when "00011110011100",
                             25654 when "00011110011101",
                             25641 when "00011110011110",
                             25628 when "00011110011111",
                             25615 when "00011110100000",
                             25602 when "00011110100001",
                             25589 when "00011110100010",
                             25575 when "00011110100011",
                             25562 when "00011110100100",
                             25549 when "00011110100101",
                             25536 when "00011110100110",
                             25523 when "00011110100111",
                             25510 when "00011110101000",
                             25497 when "00011110101001",
                             25484 when "00011110101010",
                             25471 when "00011110101011",
                             25458 when "00011110101100",
                             25445 when "00011110101101",
                             25432 when "00011110101110",
                             25419 when "00011110101111",
                             25407 when "00011110110000",
                             25394 when "00011110110001",
                             25381 when "00011110110010",
                             25368 when "00011110110011",
                             25355 when "00011110110100",
                             25342 when "00011110110101",
                             25329 when "00011110110110",
                             25316 when "00011110110111",
                             25304 when "00011110111000",
                             25291 when "00011110111001",
                             25278 when "00011110111010",
                             25265 when "00011110111011",
                             25253 when "00011110111100",
                             25240 when "00011110111101",
                             25227 when "00011110111110",
                             25214 when "00011110111111",
                             25202 when "00011111000000",
                             25189 when "00011111000001",
                             25176 when "00011111000010",
                             25164 when "00011111000011",
                             25151 when "00011111000100",
                             25138 when "00011111000101",
                             25126 when "00011111000110",
                             25113 when "00011111000111",
                             25100 when "00011111001000",
                             25088 when "00011111001001",
                             25075 when "00011111001010",
                             25063 when "00011111001011",
                             25050 when "00011111001100",
                             25038 when "00011111001101",
                             25025 when "00011111001110",
                             25013 when "00011111001111",
                             25000 when "00011111010000",
                             24988 when "00011111010001",
                             24975 when "00011111010010",
                             24963 when "00011111010011",
                             24950 when "00011111010100",
                             24938 when "00011111010101",
                             24925 when "00011111010110",
                             24913 when "00011111010111",
                             24900 when "00011111011000",
                             24888 when "00011111011001",
                             24876 when "00011111011010",
                             24863 when "00011111011011",
                             24851 when "00011111011100",
                             24839 when "00011111011101",
                             24826 when "00011111011110",
                             24814 when "00011111011111",
                             24802 when "00011111100000",
                             24789 when "00011111100001",
                             24777 when "00011111100010",
                             24765 when "00011111100011",
                             24752 when "00011111100100",
                             24740 when "00011111100101",
                             24728 when "00011111100110",
                             24716 when "00011111100111",
                             24704 when "00011111101000",
                             24691 when "00011111101001",
                             24679 when "00011111101010",
                             24667 when "00011111101011",
                             24655 when "00011111101100",
                             24643 when "00011111101101",
                             24631 when "00011111101110",
                             24618 when "00011111101111",
                             24606 when "00011111110000",
                             24594 when "00011111110001",
                             24582 when "00011111110010",
                             24570 when "00011111110011",
                             24558 when "00011111110100",
                             24546 when "00011111110101",
                             24534 when "00011111110110",
                             24522 when "00011111110111",
                             24510 when "00011111111000",
                             24498 when "00011111111001",
                             24486 when "00011111111010",
                             24474 when "00011111111011",
                             24462 when "00011111111100",
                             24450 when "00011111111101",
                             24438 when "00011111111110",
                             24426 when "00011111111111",
                             24414 when "00100000000000",
                             24402 when "00100000000001",
                             24390 when "00100000000010",
                             24378 when "00100000000011",
                             24366 when "00100000000100",
                             24355 when "00100000000101",
                             24343 when "00100000000110",
                             24331 when "00100000000111",
                             24319 when "00100000001000",
                             24307 when "00100000001001",
                             24295 when "00100000001010",
                             24284 when "00100000001011",
                             24272 when "00100000001100",
                             24260 when "00100000001101",
                             24248 when "00100000001110",
                             24237 when "00100000001111",
                             24225 when "00100000010000",
                             24213 when "00100000010001",
                             24201 when "00100000010010",
                             24190 when "00100000010011",
                             24178 when "00100000010100",
                             24166 when "00100000010101",
                             24155 when "00100000010110",
                             24143 when "00100000010111",
                             24131 when "00100000011000",
                             24120 when "00100000011001",
                             24108 when "00100000011010",
                             24096 when "00100000011011",
                             24085 when "00100000011100",
                             24073 when "00100000011101",
                             24062 when "00100000011110",
                             24050 when "00100000011111",
                             24038 when "00100000100000",
                             24027 when "00100000100001",
                             24015 when "00100000100010",
                             24004 when "00100000100011",
                             23992 when "00100000100100",
                             23981 when "00100000100101",
                             23969 when "00100000100110",
                             23958 when "00100000100111",
                             23946 when "00100000101000",
                             23935 when "00100000101001",
                             23923 when "00100000101010",
                             23912 when "00100000101011",
                             23901 when "00100000101100",
                             23889 when "00100000101101",
                             23878 when "00100000101110",
                             23866 when "00100000101111",
                             23855 when "00100000110000",
                             23844 when "00100000110001",
                             23832 when "00100000110010",
                             23821 when "00100000110011",
                             23810 when "00100000110100",
                             23798 when "00100000110101",
                             23787 when "00100000110110",
                             23776 when "00100000110111",
                             23764 when "00100000111000",
                             23753 when "00100000111001",
                             23742 when "00100000111010",
                             23730 when "00100000111011",
                             23719 when "00100000111100",
                             23708 when "00100000111101",
                             23697 when "00100000111110",
                             23685 when "00100000111111",
                             23674 when "00100001000000",
                             23663 when "00100001000001",
                             23652 when "00100001000010",
                             23641 when "00100001000011",
                             23629 when "00100001000100",
                             23618 when "00100001000101",
                             23607 when "00100001000110",
                             23596 when "00100001000111",
                             23585 when "00100001001000",
                             23574 when "00100001001001",
                             23563 when "00100001001010",
                             23552 when "00100001001011",
                             23540 when "00100001001100",
                             23529 when "00100001001101",
                             23518 when "00100001001110",
                             23507 when "00100001001111",
                             23496 when "00100001010000",
                             23485 when "00100001010001",
                             23474 when "00100001010010",
                             23463 when "00100001010011",
                             23452 when "00100001010100",
                             23441 when "00100001010101",
                             23430 when "00100001010110",
                             23419 when "00100001010111",
                             23408 when "00100001011000",
                             23397 when "00100001011001",
                             23386 when "00100001011010",
                             23375 when "00100001011011",
                             23364 when "00100001011100",
                             23354 when "00100001011101",
                             23343 when "00100001011110",
                             23332 when "00100001011111",
                             23321 when "00100001100000",
                             23310 when "00100001100001",
                             23299 when "00100001100010",
                             23288 when "00100001100011",
                             23277 when "00100001100100",
                             23267 when "00100001100101",
                             23256 when "00100001100110",
                             23245 when "00100001100111",
                             23234 when "00100001101000",
                             23223 when "00100001101001",
                             23213 when "00100001101010",
                             23202 when "00100001101011",
                             23191 when "00100001101100",
                             23180 when "00100001101101",
                             23170 when "00100001101110",
                             23159 when "00100001101111",
                             23148 when "00100001110000",
                             23137 when "00100001110001",
                             23127 when "00100001110010",
                             23116 when "00100001110011",
                             23105 when "00100001110100",
                             23095 when "00100001110101",
                             23084 when "00100001110110",
                             23073 when "00100001110111",
                             23063 when "00100001111000",
                             23052 when "00100001111001",
                             23041 when "00100001111010",
                             23031 when "00100001111011",
                             23020 when "00100001111100",
                             23010 when "00100001111101",
                             22999 when "00100001111110",
                             22989 when "00100001111111",
                             22978 when "00100010000000",
                             22967 when "00100010000001",
                             22957 when "00100010000010",
                             22946 when "00100010000011",
                             22936 when "00100010000100",
                             22925 when "00100010000101",
                             22915 when "00100010000110",
                             22904 when "00100010000111",
                             22894 when "00100010001000",
                             22883 when "00100010001001",
                             22873 when "00100010001010",
                             22862 when "00100010001011",
                             22852 when "00100010001100",
                             22841 when "00100010001101",
                             22831 when "00100010001110",
                             22821 when "00100010001111",
                             22810 when "00100010010000",
                             22800 when "00100010010001",
                             22789 when "00100010010010",
                             22779 when "00100010010011",
                             22769 when "00100010010100",
                             22758 when "00100010010101",
                             22748 when "00100010010110",
                             22738 when "00100010010111",
                             22727 when "00100010011000",
                             22717 when "00100010011001",
                             22707 when "00100010011010",
                             22696 when "00100010011011",
                             22686 when "00100010011100",
                             22676 when "00100010011101",
                             22665 when "00100010011110",
                             22655 when "00100010011111",
                             22645 when "00100010100000",
                             22635 when "00100010100001",
                             22624 when "00100010100010",
                             22614 when "00100010100011",
                             22604 when "00100010100100",
                             22594 when "00100010100101",
                             22584 when "00100010100110",
                             22573 when "00100010100111",
                             22563 when "00100010101000",
                             22553 when "00100010101001",
                             22543 when "00100010101010",
                             22533 when "00100010101011",
                             22523 when "00100010101100",
                             22512 when "00100010101101",
                             22502 when "00100010101110",
                             22492 when "00100010101111",
                             22482 when "00100010110000",
                             22472 when "00100010110001",
                             22462 when "00100010110010",
                             22452 when "00100010110011",
                             22442 when "00100010110100",
                             22432 when "00100010110101",
                             22422 when "00100010110110",
                             22411 when "00100010110111",
                             22401 when "00100010111000",
                             22391 when "00100010111001",
                             22381 when "00100010111010",
                             22371 when "00100010111011",
                             22361 when "00100010111100",
                             22351 when "00100010111101",
                             22341 when "00100010111110",
                             22331 when "00100010111111",
                             22321 when "00100011000000",
                             22311 when "00100011000001",
                             22302 when "00100011000010",
                             22292 when "00100011000011",
                             22282 when "00100011000100",
                             22272 when "00100011000101",
                             22262 when "00100011000110",
                             22252 when "00100011000111",
                             22242 when "00100011001000",
                             22232 when "00100011001001",
                             22222 when "00100011001010",
                             22212 when "00100011001011",
                             22202 when "00100011001100",
                             22193 when "00100011001101",
                             22183 when "00100011001110",
                             22173 when "00100011001111",
                             22163 when "00100011010000",
                             22153 when "00100011010001",
                             22143 when "00100011010010",
                             22134 when "00100011010011",
                             22124 when "00100011010100",
                             22114 when "00100011010101",
                             22104 when "00100011010110",
                             22095 when "00100011010111",
                             22085 when "00100011011000",
                             22075 when "00100011011001",
                             22065 when "00100011011010",
                             22056 when "00100011011011",
                             22046 when "00100011011100",
                             22036 when "00100011011101",
                             22026 when "00100011011110",
                             22017 when "00100011011111",
                             22007 when "00100011100000",
                             21997 when "00100011100001",
                             21988 when "00100011100010",
                             21978 when "00100011100011",
                             21968 when "00100011100100",
                             21959 when "00100011100101",
                             21949 when "00100011100110",
                             21939 when "00100011100111",
                             21930 when "00100011101000",
                             21920 when "00100011101001",
                             21911 when "00100011101010",
                             21901 when "00100011101011",
                             21891 when "00100011101100",
                             21882 when "00100011101101",
                             21872 when "00100011101110",
                             21863 when "00100011101111",
                             21853 when "00100011110000",
                             21844 when "00100011110001",
                             21834 when "00100011110010",
                             21825 when "00100011110011",
                             21815 when "00100011110100",
                             21805 when "00100011110101",
                             21796 when "00100011110110",
                             21786 when "00100011110111",
                             21777 when "00100011111000",
                             21768 when "00100011111001",
                             21758 when "00100011111010",
                             21749 when "00100011111011",
                             21739 when "00100011111100",
                             21730 when "00100011111101",
                             21720 when "00100011111110",
                             21711 when "00100011111111",
                             21701 when "00100100000000",
                             21692 when "00100100000001",
                             21683 when "00100100000010",
                             21673 when "00100100000011",
                             21664 when "00100100000100",
                             21654 when "00100100000101",
                             21645 when "00100100000110",
                             21636 when "00100100000111",
                             21626 when "00100100001000",
                             21617 when "00100100001001",
                             21608 when "00100100001010",
                             21598 when "00100100001011",
                             21589 when "00100100001100",
                             21580 when "00100100001101",
                             21570 when "00100100001110",
                             21561 when "00100100001111",
                             21552 when "00100100010000",
                             21542 when "00100100010001",
                             21533 when "00100100010010",
                             21524 when "00100100010011",
                             21515 when "00100100010100",
                             21505 when "00100100010101",
                             21496 when "00100100010110",
                             21487 when "00100100010111",
                             21478 when "00100100011000",
                             21468 when "00100100011001",
                             21459 when "00100100011010",
                             21450 when "00100100011011",
                             21441 when "00100100011100",
                             21432 when "00100100011101",
                             21422 when "00100100011110",
                             21413 when "00100100011111",
                             21404 when "00100100100000",
                             21395 when "00100100100001",
                             21386 when "00100100100010",
                             21377 when "00100100100011",
                             21368 when "00100100100100",
                             21358 when "00100100100101",
                             21349 when "00100100100110",
                             21340 when "00100100100111",
                             21331 when "00100100101000",
                             21322 when "00100100101001",
                             21313 when "00100100101010",
                             21304 when "00100100101011",
                             21295 when "00100100101100",
                             21286 when "00100100101101",
                             21277 when "00100100101110",
                             21268 when "00100100101111",
                             21259 when "00100100110000",
                             21249 when "00100100110001",
                             21240 when "00100100110010",
                             21231 when "00100100110011",
                             21222 when "00100100110100",
                             21213 when "00100100110101",
                             21204 when "00100100110110",
                             21195 when "00100100110111",
                             21186 when "00100100111000",
                             21177 when "00100100111001",
                             21169 when "00100100111010",
                             21160 when "00100100111011",
                             21151 when "00100100111100",
                             21142 when "00100100111101",
                             21133 when "00100100111110",
                             21124 when "00100100111111",
                             21115 when "00100101000000",
                             21106 when "00100101000001",
                             21097 when "00100101000010",
                             21088 when "00100101000011",
                             21079 when "00100101000100",
                             21070 when "00100101000101",
                             21061 when "00100101000110",
                             21053 when "00100101000111",
                             21044 when "00100101001000",
                             21035 when "00100101001001",
                             21026 when "00100101001010",
                             21017 when "00100101001011",
                             21008 when "00100101001100",
                             21000 when "00100101001101",
                             20991 when "00100101001110",
                             20982 when "00100101001111",
                             20973 when "00100101010000",
                             20964 when "00100101010001",
                             20956 when "00100101010010",
                             20947 when "00100101010011",
                             20938 when "00100101010100",
                             20929 when "00100101010101",
                             20921 when "00100101010110",
                             20912 when "00100101010111",
                             20903 when "00100101011000",
                             20894 when "00100101011001",
                             20886 when "00100101011010",
                             20877 when "00100101011011",
                             20868 when "00100101011100",
                             20859 when "00100101011101",
                             20851 when "00100101011110",
                             20842 when "00100101011111",
                             20833 when "00100101100000",
                             20825 when "00100101100001",
                             20816 when "00100101100010",
                             20807 when "00100101100011",
                             20799 when "00100101100100",
                             20790 when "00100101100101",
                             20781 when "00100101100110",
                             20773 when "00100101100111",
                             20764 when "00100101101000",
                             20756 when "00100101101001",
                             20747 when "00100101101010",
                             20738 when "00100101101011",
                             20730 when "00100101101100",
                             20721 when "00100101101101",
                             20713 when "00100101101110",
                             20704 when "00100101101111",
                             20695 when "00100101110000",
                             20687 when "00100101110001",
                             20678 when "00100101110010",
                             20670 when "00100101110011",
                             20661 when "00100101110100",
                             20653 when "00100101110101",
                             20644 when "00100101110110",
                             20636 when "00100101110111",
                             20627 when "00100101111000",
                             20619 when "00100101111001",
                             20610 when "00100101111010",
                             20602 when "00100101111011",
                             20593 when "00100101111100",
                             20585 when "00100101111101",
                             20576 when "00100101111110",
                             20568 when "00100101111111",
                             20559 when "00100110000000",
                             20551 when "00100110000001",
                             20542 when "00100110000010",
                             20534 when "00100110000011",
                             20525 when "00100110000100",
                             20517 when "00100110000101",
                             20509 when "00100110000110",
                             20500 when "00100110000111",
                             20492 when "00100110001000",
                             20483 when "00100110001001",
                             20475 when "00100110001010",
                             20467 when "00100110001011",
                             20458 when "00100110001100",
                             20450 when "00100110001101",
                             20442 when "00100110001110",
                             20433 when "00100110001111",
                             20425 when "00100110010000",
                             20416 when "00100110010001",
                             20408 when "00100110010010",
                             20400 when "00100110010011",
                             20392 when "00100110010100",
                             20383 when "00100110010101",
                             20375 when "00100110010110",
                             20367 when "00100110010111",
                             20358 when "00100110011000",
                             20350 when "00100110011001",
                             20342 when "00100110011010",
                             20333 when "00100110011011",
                             20325 when "00100110011100",
                             20317 when "00100110011101",
                             20309 when "00100110011110",
                             20300 when "00100110011111",
                             20292 when "00100110100000",
                             20284 when "00100110100001",
                             20276 when "00100110100010",
                             20268 when "00100110100011",
                             20259 when "00100110100100",
                             20251 when "00100110100101",
                             20243 when "00100110100110",
                             20235 when "00100110100111",
                             20227 when "00100110101000",
                             20218 when "00100110101001",
                             20210 when "00100110101010",
                             20202 when "00100110101011",
                             20194 when "00100110101100",
                             20186 when "00100110101101",
                             20178 when "00100110101110",
                             20169 when "00100110101111",
                             20161 when "00100110110000",
                             20153 when "00100110110001",
                             20145 when "00100110110010",
                             20137 when "00100110110011",
                             20129 when "00100110110100",
                             20121 when "00100110110101",
                             20113 when "00100110110110",
                             20105 when "00100110110111",
                             20096 when "00100110111000",
                             20088 when "00100110111001",
                             20080 when "00100110111010",
                             20072 when "00100110111011",
                             20064 when "00100110111100",
                             20056 when "00100110111101",
                             20048 when "00100110111110",
                             20040 when "00100110111111",
                             20032 when "00100111000000",
                             20024 when "00100111000001",
                             20016 when "00100111000010",
                             20008 when "00100111000011",
                             20000 when "00100111000100",
                             19992 when "00100111000101",
                             19984 when "00100111000110",
                             19976 when "00100111000111",
                             19968 when "00100111001000",
                             19960 when "00100111001001",
                             19952 when "00100111001010",
                             19944 when "00100111001011",
                             19936 when "00100111001100",
                             19928 when "00100111001101",
                             19920 when "00100111001110",
                             19912 when "00100111001111",
                             19904 when "00100111010000",
                             19897 when "00100111010001",
                             19889 when "00100111010010",
                             19881 when "00100111010011",
                             19873 when "00100111010100",
                             19865 when "00100111010101",
                             19857 when "00100111010110",
                             19849 when "00100111010111",
                             19841 when "00100111011000",
                             19833 when "00100111011001",
                             19826 when "00100111011010",
                             19818 when "00100111011011",
                             19810 when "00100111011100",
                             19802 when "00100111011101",
                             19794 when "00100111011110",
                             19786 when "00100111011111",
                             19778 when "00100111100000",
                             19771 when "00100111100001",
                             19763 when "00100111100010",
                             19755 when "00100111100011",
                             19747 when "00100111100100",
                             19739 when "00100111100101",
                             19732 when "00100111100110",
                             19724 when "00100111100111",
                             19716 when "00100111101000",
                             19708 when "00100111101001",
                             19701 when "00100111101010",
                             19693 when "00100111101011",
                             19685 when "00100111101100",
                             19677 when "00100111101101",
                             19670 when "00100111101110",
                             19662 when "00100111101111",
                             19654 when "00100111110000",
                             19646 when "00100111110001",
                             19639 when "00100111110010",
                             19631 when "00100111110011",
                             19623 when "00100111110100",
                             19616 when "00100111110101",
                             19608 when "00100111110110",
                             19600 when "00100111110111",
                             19592 when "00100111111000",
                             19585 when "00100111111001",
                             19577 when "00100111111010",
                             19569 when "00100111111011",
                             19562 when "00100111111100",
                             19554 when "00100111111101",
                             19547 when "00100111111110",
                             19539 when "00100111111111",
                             19531 when "00101000000000",
                             19524 when "00101000000001",
                             19516 when "00101000000010",
                             19508 when "00101000000011",
                             19501 when "00101000000100",
                             19493 when "00101000000101",
                             19486 when "00101000000110",
                             19478 when "00101000000111",
                             19470 when "00101000001000",
                             19463 when "00101000001001",
                             19455 when "00101000001010",
                             19448 when "00101000001011",
                             19440 when "00101000001100",
                             19433 when "00101000001101",
                             19425 when "00101000001110",
                             19417 when "00101000001111",
                             19410 when "00101000010000",
                             19402 when "00101000010001",
                             19395 when "00101000010010",
                             19387 when "00101000010011",
                             19380 when "00101000010100",
                             19372 when "00101000010101",
                             19365 when "00101000010110",
                             19357 when "00101000010111",
                             19350 when "00101000011000",
                             19342 when "00101000011001",
                             19335 when "00101000011010",
                             19327 when "00101000011011",
                             19320 when "00101000011100",
                             19312 when "00101000011101",
                             19305 when "00101000011110",
                             19298 when "00101000011111",
                             19290 when "00101000100000",
                             19283 when "00101000100001",
                             19275 when "00101000100010",
                             19268 when "00101000100011",
                             19260 when "00101000100100",
                             19253 when "00101000100101",
                             19246 when "00101000100110",
                             19238 when "00101000100111",
                             19231 when "00101000101000",
                             19223 when "00101000101001",
                             19216 when "00101000101010",
                             19209 when "00101000101011",
                             19201 when "00101000101100",
                             19194 when "00101000101101",
                             19186 when "00101000101110",
                             19179 when "00101000101111",
                             19172 when "00101000110000",
                             19164 when "00101000110001",
                             19157 when "00101000110010",
                             19150 when "00101000110011",
                             19142 when "00101000110100",
                             19135 when "00101000110101",
                             19128 when "00101000110110",
                             19120 when "00101000110111",
                             19113 when "00101000111000",
                             19106 when "00101000111001",
                             19099 when "00101000111010",
                             19091 when "00101000111011",
                             19084 when "00101000111100",
                             19077 when "00101000111101",
                             19069 when "00101000111110",
                             19062 when "00101000111111",
                             19055 when "00101001000000",
                             19048 when "00101001000001",
                             19040 when "00101001000010",
                             19033 when "00101001000011",
                             19026 when "00101001000100",
                             19019 when "00101001000101",
                             19011 when "00101001000110",
                             19004 when "00101001000111",
                             18997 when "00101001001000",
                             18990 when "00101001001001",
                             18983 when "00101001001010",
                             18975 when "00101001001011",
                             18968 when "00101001001100",
                             18961 when "00101001001101",
                             18954 when "00101001001110",
                             18947 when "00101001001111",
                             18939 when "00101001010000",
                             18932 when "00101001010001",
                             18925 when "00101001010010",
                             18918 when "00101001010011",
                             18911 when "00101001010100",
                             18904 when "00101001010101",
                             18896 when "00101001010110",
                             18889 when "00101001010111",
                             18882 when "00101001011000",
                             18875 when "00101001011001",
                             18868 when "00101001011010",
                             18861 when "00101001011011",
                             18854 when "00101001011100",
                             18847 when "00101001011101",
                             18839 when "00101001011110",
                             18832 when "00101001011111",
                             18825 when "00101001100000",
                             18818 when "00101001100001",
                             18811 when "00101001100010",
                             18804 when "00101001100011",
                             18797 when "00101001100100",
                             18790 when "00101001100101",
                             18783 when "00101001100110",
                             18776 when "00101001100111",
                             18769 when "00101001101000",
                             18762 when "00101001101001",
                             18755 when "00101001101010",
                             18748 when "00101001101011",
                             18741 when "00101001101100",
                             18734 when "00101001101101",
                             18727 when "00101001101110",
                             18720 when "00101001101111",
                             18713 when "00101001110000",
                             18706 when "00101001110001",
                             18699 when "00101001110010",
                             18692 when "00101001110011",
                             18685 when "00101001110100",
                             18678 when "00101001110101",
                             18671 when "00101001110110",
                             18664 when "00101001110111",
                             18657 when "00101001111000",
                             18650 when "00101001111001",
                             18643 when "00101001111010",
                             18636 when "00101001111011",
                             18629 when "00101001111100",
                             18622 when "00101001111101",
                             18615 when "00101001111110",
                             18608 when "00101001111111",
                             18601 when "00101010000000",
                             18594 when "00101010000001",
                             18587 when "00101010000010",
                             18580 when "00101010000011",
                             18574 when "00101010000100",
                             18567 when "00101010000101",
                             18560 when "00101010000110",
                             18553 when "00101010000111",
                             18546 when "00101010001000",
                             18539 when "00101010001001",
                             18532 when "00101010001010",
                             18525 when "00101010001011",
                             18519 when "00101010001100",
                             18512 when "00101010001101",
                             18505 when "00101010001110",
                             18498 when "00101010001111",
                             18491 when "00101010010000",
                             18484 when "00101010010001",
                             18477 when "00101010010010",
                             18471 when "00101010010011",
                             18464 when "00101010010100",
                             18457 when "00101010010101",
                             18450 when "00101010010110",
                             18443 when "00101010010111",
                             18437 when "00101010011000",
                             18430 when "00101010011001",
                             18423 when "00101010011010",
                             18416 when "00101010011011",
                             18409 when "00101010011100",
                             18403 when "00101010011101",
                             18396 when "00101010011110",
                             18389 when "00101010011111",
                             18382 when "00101010100000",
                             18376 when "00101010100001",
                             18369 when "00101010100010",
                             18362 when "00101010100011",
                             18355 when "00101010100100",
                             18349 when "00101010100101",
                             18342 when "00101010100110",
                             18335 when "00101010100111",
                             18328 when "00101010101000",
                             18322 when "00101010101001",
                             18315 when "00101010101010",
                             18308 when "00101010101011",
                             18302 when "00101010101100",
                             18295 when "00101010101101",
                             18288 when "00101010101110",
                             18282 when "00101010101111",
                             18275 when "00101010110000",
                             18268 when "00101010110001",
                             18262 when "00101010110010",
                             18255 when "00101010110011",
                             18248 when "00101010110100",
                             18242 when "00101010110101",
                             18235 when "00101010110110",
                             18228 when "00101010110111",
                             18222 when "00101010111000",
                             18215 when "00101010111001",
                             18208 when "00101010111010",
                             18202 when "00101010111011",
                             18195 when "00101010111100",
                             18188 when "00101010111101",
                             18182 when "00101010111110",
                             18175 when "00101010111111",
                             18169 when "00101011000000",
                             18162 when "00101011000001",
                             18155 when "00101011000010",
                             18149 when "00101011000011",
                             18142 when "00101011000100",
                             18136 when "00101011000101",
                             18129 when "00101011000110",
                             18123 when "00101011000111",
                             18116 when "00101011001000",
                             18109 when "00101011001001",
                             18103 when "00101011001010",
                             18096 when "00101011001011",
                             18090 when "00101011001100",
                             18083 when "00101011001101",
                             18077 when "00101011001110",
                             18070 when "00101011001111",
                             18064 when "00101011010000",
                             18057 when "00101011010001",
                             18051 when "00101011010010",
                             18044 when "00101011010011",
                             18038 when "00101011010100",
                             18031 when "00101011010101",
                             18025 when "00101011010110",
                             18018 when "00101011010111",
                             18012 when "00101011011000",
                             18005 when "00101011011001",
                             17999 when "00101011011010",
                             17992 when "00101011011011",
                             17986 when "00101011011100",
                             17979 when "00101011011101",
                             17973 when "00101011011110",
                             17966 when "00101011011111",
                             17960 when "00101011100000",
                             17953 when "00101011100001",
                             17947 when "00101011100010",
                             17940 when "00101011100011",
                             17934 when "00101011100100",
                             17928 when "00101011100101",
                             17921 when "00101011100110",
                             17915 when "00101011100111",
                             17908 when "00101011101000",
                             17902 when "00101011101001",
                             17895 when "00101011101010",
                             17889 when "00101011101011",
                             17883 when "00101011101100",
                             17876 when "00101011101101",
                             17870 when "00101011101110",
                             17864 when "00101011101111",
                             17857 when "00101011110000",
                             17851 when "00101011110001",
                             17844 when "00101011110010",
                             17838 when "00101011110011",
                             17832 when "00101011110100",
                             17825 when "00101011110101",
                             17819 when "00101011110110",
                             17813 when "00101011110111",
                             17806 when "00101011111000",
                             17800 when "00101011111001",
                             17794 when "00101011111010",
                             17787 when "00101011111011",
                             17781 when "00101011111100",
                             17775 when "00101011111101",
                             17768 when "00101011111110",
                             17762 when "00101011111111",
                             17756 when "00101100000000",
                             17749 when "00101100000001",
                             17743 when "00101100000010",
                             17737 when "00101100000011",
                             17730 when "00101100000100",
                             17724 when "00101100000101",
                             17718 when "00101100000110",
                             17712 when "00101100000111",
                             17705 when "00101100001000",
                             17699 when "00101100001001",
                             17693 when "00101100001010",
                             17687 when "00101100001011",
                             17680 when "00101100001100",
                             17674 when "00101100001101",
                             17668 when "00101100001110",
                             17662 when "00101100001111",
                             17655 when "00101100010000",
                             17649 when "00101100010001",
                             17643 when "00101100010010",
                             17637 when "00101100010011",
                             17630 when "00101100010100",
                             17624 when "00101100010101",
                             17618 when "00101100010110",
                             17612 when "00101100010111",
                             17606 when "00101100011000",
                             17599 when "00101100011001",
                             17593 when "00101100011010",
                             17587 when "00101100011011",
                             17581 when "00101100011100",
                             17575 when "00101100011101",
                             17569 when "00101100011110",
                             17562 when "00101100011111",
                             17556 when "00101100100000",
                             17550 when "00101100100001",
                             17544 when "00101100100010",
                             17538 when "00101100100011",
                             17532 when "00101100100100",
                             17525 when "00101100100101",
                             17519 when "00101100100110",
                             17513 when "00101100100111",
                             17507 when "00101100101000",
                             17501 when "00101100101001",
                             17495 when "00101100101010",
                             17489 when "00101100101011",
                             17483 when "00101100101100",
                             17476 when "00101100101101",
                             17470 when "00101100101110",
                             17464 when "00101100101111",
                             17458 when "00101100110000",
                             17452 when "00101100110001",
                             17446 when "00101100110010",
                             17440 when "00101100110011",
                             17434 when "00101100110100",
                             17428 when "00101100110101",
                             17422 when "00101100110110",
                             17416 when "00101100110111",
                             17409 when "00101100111000",
                             17403 when "00101100111001",
                             17397 when "00101100111010",
                             17391 when "00101100111011",
                             17385 when "00101100111100",
                             17379 when "00101100111101",
                             17373 when "00101100111110",
                             17367 when "00101100111111",
                             17361 when "00101101000000",
                             17355 when "00101101000001",
                             17349 when "00101101000010",
                             17343 when "00101101000011",
                             17337 when "00101101000100",
                             17331 when "00101101000101",
                             17325 when "00101101000110",
                             17319 when "00101101000111",
                             17313 when "00101101001000",
                             17307 when "00101101001001",
                             17301 when "00101101001010",
                             17295 when "00101101001011",
                             17289 when "00101101001100",
                             17283 when "00101101001101",
                             17277 when "00101101001110",
                             17271 when "00101101001111",
                             17265 when "00101101010000",
                             17259 when "00101101010001",
                             17253 when "00101101010010",
                             17247 when "00101101010011",
                             17241 when "00101101010100",
                             17235 when "00101101010101",
                             17229 when "00101101010110",
                             17224 when "00101101010111",
                             17218 when "00101101011000",
                             17212 when "00101101011001",
                             17206 when "00101101011010",
                             17200 when "00101101011011",
                             17194 when "00101101011100",
                             17188 when "00101101011101",
                             17182 when "00101101011110",
                             17176 when "00101101011111",
                             17170 when "00101101100000",
                             17164 when "00101101100001",
                             17159 when "00101101100010",
                             17153 when "00101101100011",
                             17147 when "00101101100100",
                             17141 when "00101101100101",
                             17135 when "00101101100110",
                             17129 when "00101101100111",
                             17123 when "00101101101000",
                             17117 when "00101101101001",
                             17112 when "00101101101010",
                             17106 when "00101101101011",
                             17100 when "00101101101100",
                             17094 when "00101101101101",
                             17088 when "00101101101110",
                             17082 when "00101101101111",
                             17077 when "00101101110000",
                             17071 when "00101101110001",
                             17065 when "00101101110010",
                             17059 when "00101101110011",
                             17053 when "00101101110100",
                             17047 when "00101101110101",
                             17042 when "00101101110110",
                             17036 when "00101101110111",
                             17030 when "00101101111000",
                             17024 when "00101101111001",
                             17018 when "00101101111010",
                             17013 when "00101101111011",
                             17007 when "00101101111100",
                             17001 when "00101101111101",
                             16995 when "00101101111110",
                             16989 when "00101101111111",
                             16984 when "00101110000000",
                             16978 when "00101110000001",
                             16972 when "00101110000010",
                             16966 when "00101110000011",
                             16961 when "00101110000100",
                             16955 when "00101110000101",
                             16949 when "00101110000110",
                             16943 when "00101110000111",
                             16938 when "00101110001000",
                             16932 when "00101110001001",
                             16926 when "00101110001010",
                             16920 when "00101110001011",
                             16915 when "00101110001100",
                             16909 when "00101110001101",
                             16903 when "00101110001110",
                             16898 when "00101110001111",
                             16892 when "00101110010000",
                             16886 when "00101110010001",
                             16880 when "00101110010010",
                             16875 when "00101110010011",
                             16869 when "00101110010100",
                             16863 when "00101110010101",
                             16858 when "00101110010110",
                             16852 when "00101110010111",
                             16846 when "00101110011000",
                             16841 when "00101110011001",
                             16835 when "00101110011010",
                             16829 when "00101110011011",
                             16824 when "00101110011100",
                             16818 when "00101110011101",
                             16812 when "00101110011110",
                             16807 when "00101110011111",
                             16801 when "00101110100000",
                             16795 when "00101110100001",
                             16790 when "00101110100010",
                             16784 when "00101110100011",
                             16779 when "00101110100100",
                             16773 when "00101110100101",
                             16767 when "00101110100110",
                             16762 when "00101110100111",
                             16756 when "00101110101000",
                             16750 when "00101110101001",
                             16745 when "00101110101010",
                             16739 when "00101110101011",
                             16734 when "00101110101100",
                             16728 when "00101110101101",
                             16722 when "00101110101110",
                             16717 when "00101110101111",
                             16711 when "00101110110000",
                             16706 when "00101110110001",
                             16700 when "00101110110010",
                             16694 when "00101110110011",
                             16689 when "00101110110100",
                             16683 when "00101110110101",
                             16678 when "00101110110110",
                             16672 when "00101110110111",
                             16667 when "00101110111000",
                             16661 when "00101110111001",
                             16656 when "00101110111010",
                             16650 when "00101110111011",
                             16644 when "00101110111100",
                             16639 when "00101110111101",
                             16633 when "00101110111110",
                             16628 when "00101110111111",
                             16622 when "00101111000000",
                             16617 when "00101111000001",
                             16611 when "00101111000010",
                             16606 when "00101111000011",
                             16600 when "00101111000100",
                             16595 when "00101111000101",
                             16589 when "00101111000110",
                             16584 when "00101111000111",
                             16578 when "00101111001000",
                             16573 when "00101111001001",
                             16567 when "00101111001010",
                             16562 when "00101111001011",
                             16556 when "00101111001100",
                             16551 when "00101111001101",
                             16545 when "00101111001110",
                             16540 when "00101111001111",
                             16534 when "00101111010000",
                             16529 when "00101111010001",
                             16523 when "00101111010010",
                             16518 when "00101111010011",
                             16513 when "00101111010100",
                             16507 when "00101111010101",
                             16502 when "00101111010110",
                             16496 when "00101111010111",
                             16491 when "00101111011000",
                             16485 when "00101111011001",
                             16480 when "00101111011010",
                             16474 when "00101111011011",
                             16469 when "00101111011100",
                             16464 when "00101111011101",
                             16458 when "00101111011110",
                             16453 when "00101111011111",
                             16447 when "00101111100000",
                             16442 when "00101111100001",
                             16437 when "00101111100010",
                             16431 when "00101111100011",
                             16426 when "00101111100100",
                             16420 when "00101111100101",
                             16415 when "00101111100110",
                             16410 when "00101111100111",
                             16404 when "00101111101000",
                             16399 when "00101111101001",
                             16393 when "00101111101010",
                             16388 when "00101111101011",
                             16383 when "00101111101100",
                             16377 when "00101111101101",
                             16372 when "00101111101110",
                             16367 when "00101111101111",
                             16361 when "00101111110000",
                             16356 when "00101111110001",
                             16351 when "00101111110010",
                             16345 when "00101111110011",
                             16340 when "00101111110100",
                             16335 when "00101111110101",
                             16329 when "00101111110110",
                             16324 when "00101111110111",
                             16319 when "00101111111000",
                             16313 when "00101111111001",
                             16308 when "00101111111010",
                             16303 when "00101111111011",
                             16297 when "00101111111100",
                             16292 when "00101111111101",
                             16287 when "00101111111110",
                             16281 when "00101111111111",
                             16276 when "00110000000000",
                             16271 when "00110000000001",
                             16265 when "00110000000010",
                             16260 when "00110000000011",
                             16255 when "00110000000100",
                             16250 when "00110000000101",
                             16244 when "00110000000110",
                             16239 when "00110000000111",
                             16234 when "00110000001000",
                             16228 when "00110000001001",
                             16223 when "00110000001010",
                             16218 when "00110000001011",
                             16213 when "00110000001100",
                             16207 when "00110000001101",
                             16202 when "00110000001110",
                             16197 when "00110000001111",
                             16192 when "00110000010000",
                             16186 when "00110000010001",
                             16181 when "00110000010010",
                             16176 when "00110000010011",
                             16171 when "00110000010100",
                             16166 when "00110000010101",
                             16160 when "00110000010110",
                             16155 when "00110000010111",
                             16150 when "00110000011000",
                             16145 when "00110000011001",
                             16139 when "00110000011010",
                             16134 when "00110000011011",
                             16129 when "00110000011100",
                             16124 when "00110000011101",
                             16119 when "00110000011110",
                             16113 when "00110000011111",
                             16108 when "00110000100000",
                             16103 when "00110000100001",
                             16098 when "00110000100010",
                             16093 when "00110000100011",
                             16088 when "00110000100100",
                             16082 when "00110000100101",
                             16077 when "00110000100110",
                             16072 when "00110000100111",
                             16067 when "00110000101000",
                             16062 when "00110000101001",
                             16057 when "00110000101010",
                             16051 when "00110000101011",
                             16046 when "00110000101100",
                             16041 when "00110000101101",
                             16036 when "00110000101110",
                             16031 when "00110000101111",
                             16026 when "00110000110000",
                             16021 when "00110000110001",
                             16015 when "00110000110010",
                             16010 when "00110000110011",
                             16005 when "00110000110100",
                             16000 when "00110000110101",
                             15995 when "00110000110110",
                             15990 when "00110000110111",
                             15985 when "00110000111000",
                             15980 when "00110000111001",
                             15974 when "00110000111010",
                             15969 when "00110000111011",
                             15964 when "00110000111100",
                             15959 when "00110000111101",
                             15954 when "00110000111110",
                             15949 when "00110000111111",
                             15944 when "00110001000000",
                             15939 when "00110001000001",
                             15934 when "00110001000010",
                             15929 when "00110001000011",
                             15924 when "00110001000100",
                             15918 when "00110001000101",
                             15913 when "00110001000110",
                             15908 when "00110001000111",
                             15903 when "00110001001000",
                             15898 when "00110001001001",
                             15893 when "00110001001010",
                             15888 when "00110001001011",
                             15883 when "00110001001100",
                             15878 when "00110001001101",
                             15873 when "00110001001110",
                             15868 when "00110001001111",
                             15863 when "00110001010000",
                             15858 when "00110001010001",
                             15853 when "00110001010010",
                             15848 when "00110001010011",
                             15843 when "00110001010100",
                             15838 when "00110001010101",
                             15833 when "00110001010110",
                             15828 when "00110001010111",
                             15823 when "00110001011000",
                             15818 when "00110001011001",
                             15813 when "00110001011010",
                             15808 when "00110001011011",
                             15803 when "00110001011100",
                             15798 when "00110001011101",
                             15793 when "00110001011110",
                             15788 when "00110001011111",
                             15783 when "00110001100000",
                             15778 when "00110001100001",
                             15773 when "00110001100010",
                             15768 when "00110001100011",
                             15763 when "00110001100100",
                             15758 when "00110001100101",
                             15753 when "00110001100110",
                             15748 when "00110001100111",
                             15743 when "00110001101000",
                             15738 when "00110001101001",
                             15733 when "00110001101010",
                             15728 when "00110001101011",
                             15723 when "00110001101100",
                             15718 when "00110001101101",
                             15713 when "00110001101110",
                             15708 when "00110001101111",
                             15704 when "00110001110000",
                             15699 when "00110001110001",
                             15694 when "00110001110010",
                             15689 when "00110001110011",
                             15684 when "00110001110100",
                             15679 when "00110001110101",
                             15674 when "00110001110110",
                             15669 when "00110001110111",
                             15664 when "00110001111000",
                             15659 when "00110001111001",
                             15654 when "00110001111010",
                             15649 when "00110001111011",
                             15645 when "00110001111100",
                             15640 when "00110001111101",
                             15635 when "00110001111110",
                             15630 when "00110001111111",
                             15625 when "00110010000000",
                             15620 when "00110010000001",
                             15615 when "00110010000010",
                             15610 when "00110010000011",
                             15605 when "00110010000100",
                             15601 when "00110010000101",
                             15596 when "00110010000110",
                             15591 when "00110010000111",
                             15586 when "00110010001000",
                             15581 when "00110010001001",
                             15576 when "00110010001010",
                             15571 when "00110010001011",
                             15567 when "00110010001100",
                             15562 when "00110010001101",
                             15557 when "00110010001110",
                             15552 when "00110010001111",
                             15547 when "00110010010000",
                             15542 when "00110010010001",
                             15538 when "00110010010010",
                             15533 when "00110010010011",
                             15528 when "00110010010100",
                             15523 when "00110010010101",
                             15518 when "00110010010110",
                             15513 when "00110010010111",
                             15509 when "00110010011000",
                             15504 when "00110010011001",
                             15499 when "00110010011010",
                             15494 when "00110010011011",
                             15489 when "00110010011100",
                             15485 when "00110010011101",
                             15480 when "00110010011110",
                             15475 when "00110010011111",
                             15470 when "00110010100000",
                             15466 when "00110010100001",
                             15461 when "00110010100010",
                             15456 when "00110010100011",
                             15451 when "00110010100100",
                             15446 when "00110010100101",
                             15442 when "00110010100110",
                             15437 when "00110010100111",
                             15432 when "00110010101000",
                             15427 when "00110010101001",
                             15423 when "00110010101010",
                             15418 when "00110010101011",
                             15413 when "00110010101100",
                             15408 when "00110010101101",
                             15404 when "00110010101110",
                             15399 when "00110010101111",
                             15394 when "00110010110000",
                             15389 when "00110010110001",
                             15385 when "00110010110010",
                             15380 when "00110010110011",
                             15375 when "00110010110100",
                             15370 when "00110010110101",
                             15366 when "00110010110110",
                             15361 when "00110010110111",
                             15356 when "00110010111000",
                             15352 when "00110010111001",
                             15347 when "00110010111010",
                             15342 when "00110010111011",
                             15337 when "00110010111100",
                             15333 when "00110010111101",
                             15328 when "00110010111110",
                             15323 when "00110010111111",
                             15319 when "00110011000000",
                             15314 when "00110011000001",
                             15309 when "00110011000010",
                             15305 when "00110011000011",
                             15300 when "00110011000100",
                             15295 when "00110011000101",
                             15291 when "00110011000110",
                             15286 when "00110011000111",
                             15281 when "00110011001000",
                             15277 when "00110011001001",
                             15272 when "00110011001010",
                             15267 when "00110011001011",
                             15263 when "00110011001100",
                             15258 when "00110011001101",
                             15253 when "00110011001110",
                             15249 when "00110011001111",
                             15244 when "00110011010000",
                             15239 when "00110011010001",
                             15235 when "00110011010010",
                             15230 when "00110011010011",
                             15225 when "00110011010100",
                             15221 when "00110011010101",
                             15216 when "00110011010110",
                             15211 when "00110011010111",
                             15207 when "00110011011000",
                             15202 when "00110011011001",
                             15198 when "00110011011010",
                             15193 when "00110011011011",
                             15188 when "00110011011100",
                             15184 when "00110011011101",
                             15179 when "00110011011110",
                             15175 when "00110011011111",
                             15170 when "00110011100000",
                             15165 when "00110011100001",
                             15161 when "00110011100010",
                             15156 when "00110011100011",
                             15152 when "00110011100100",
                             15147 when "00110011100101",
                             15142 when "00110011100110",
                             15138 when "00110011100111",
                             15133 when "00110011101000",
                             15129 when "00110011101001",
                             15124 when "00110011101010",
                             15119 when "00110011101011",
                             15115 when "00110011101100",
                             15110 when "00110011101101",
                             15106 when "00110011101110",
                             15101 when "00110011101111",
                             15097 when "00110011110000",
                             15092 when "00110011110001",
                             15088 when "00110011110010",
                             15083 when "00110011110011",
                             15078 when "00110011110100",
                             15074 when "00110011110101",
                             15069 when "00110011110110",
                             15065 when "00110011110111",
                             15060 when "00110011111000",
                             15056 when "00110011111001",
                             15051 when "00110011111010",
                             15047 when "00110011111011",
                             15042 when "00110011111100",
                             15038 when "00110011111101",
                             15033 when "00110011111110",
                             15029 when "00110011111111",
                             15024 when "00110100000000",
                             15020 when "00110100000001",
                             15015 when "00110100000010",
                             15011 when "00110100000011",
                             15006 when "00110100000100",
                             15002 when "00110100000101",
                             14997 when "00110100000110",
                             14993 when "00110100000111",
                             14988 when "00110100001000",
                             14984 when "00110100001001",
                             14979 when "00110100001010",
                             14975 when "00110100001011",
                             14970 when "00110100001100",
                             14966 when "00110100001101",
                             14961 when "00110100001110",
                             14957 when "00110100001111",
                             14952 when "00110100010000",
                             14948 when "00110100010001",
                             14943 when "00110100010010",
                             14939 when "00110100010011",
                             14934 when "00110100010100",
                             14930 when "00110100010101",
                             14925 when "00110100010110",
                             14921 when "00110100010111",
                             14916 when "00110100011000",
                             14912 when "00110100011001",
                             14908 when "00110100011010",
                             14903 when "00110100011011",
                             14899 when "00110100011100",
                             14894 when "00110100011101",
                             14890 when "00110100011110",
                             14885 when "00110100011111",
                             14881 when "00110100100000",
                             14877 when "00110100100001",
                             14872 when "00110100100010",
                             14868 when "00110100100011",
                             14863 when "00110100100100",
                             14859 when "00110100100101",
                             14854 when "00110100100110",
                             14850 when "00110100100111",
                             14846 when "00110100101000",
                             14841 when "00110100101001",
                             14837 when "00110100101010",
                             14832 when "00110100101011",
                             14828 when "00110100101100",
                             14824 when "00110100101101",
                             14819 when "00110100101110",
                             14815 when "00110100101111",
                             14810 when "00110100110000",
                             14806 when "00110100110001",
                             14802 when "00110100110010",
                             14797 when "00110100110011",
                             14793 when "00110100110100",
                             14789 when "00110100110101",
                             14784 when "00110100110110",
                             14780 when "00110100110111",
                             14775 when "00110100111000",
                             14771 when "00110100111001",
                             14767 when "00110100111010",
                             14762 when "00110100111011",
                             14758 when "00110100111100",
                             14754 when "00110100111101",
                             14749 when "00110100111110",
                             14745 when "00110100111111",
                             14741 when "00110101000000",
                             14736 when "00110101000001",
                             14732 when "00110101000010",
                             14728 when "00110101000011",
                             14723 when "00110101000100",
                             14719 when "00110101000101",
                             14715 when "00110101000110",
                             14710 when "00110101000111",
                             14706 when "00110101001000",
                             14702 when "00110101001001",
                             14697 when "00110101001010",
                             14693 when "00110101001011",
                             14689 when "00110101001100",
                             14684 when "00110101001101",
                             14680 when "00110101001110",
                             14676 when "00110101001111",
                             14671 when "00110101010000",
                             14667 when "00110101010001",
                             14663 when "00110101010010",
                             14658 when "00110101010011",
                             14654 when "00110101010100",
                             14650 when "00110101010101",
                             14646 when "00110101010110",
                             14641 when "00110101010111",
                             14637 when "00110101011000",
                             14633 when "00110101011001",
                             14628 when "00110101011010",
                             14624 when "00110101011011",
                             14620 when "00110101011100",
                             14616 when "00110101011101",
                             14611 when "00110101011110",
                             14607 when "00110101011111",
                             14603 when "00110101100000",
                             14599 when "00110101100001",
                             14594 when "00110101100010",
                             14590 when "00110101100011",
                             14586 when "00110101100100",
                             14582 when "00110101100101",
                             14577 when "00110101100110",
                             14573 when "00110101100111",
                             14569 when "00110101101000",
                             14565 when "00110101101001",
                             14560 when "00110101101010",
                             14556 when "00110101101011",
                             14552 when "00110101101100",
                             14548 when "00110101101101",
                             14543 when "00110101101110",
                             14539 when "00110101101111",
                             14535 when "00110101110000",
                             14531 when "00110101110001",
                             14526 when "00110101110010",
                             14522 when "00110101110011",
                             14518 when "00110101110100",
                             14514 when "00110101110101",
                             14510 when "00110101110110",
                             14505 when "00110101110111",
                             14501 when "00110101111000",
                             14497 when "00110101111001",
                             14493 when "00110101111010",
                             14489 when "00110101111011",
                             14484 when "00110101111100",
                             14480 when "00110101111101",
                             14476 when "00110101111110",
                             14472 when "00110101111111",
                             14468 when "00110110000000",
                             14463 when "00110110000001",
                             14459 when "00110110000010",
                             14455 when "00110110000011",
                             14451 when "00110110000100",
                             14447 when "00110110000101",
                             14443 when "00110110000110",
                             14438 when "00110110000111",
                             14434 when "00110110001000",
                             14430 when "00110110001001",
                             14426 when "00110110001010",
                             14422 when "00110110001011",
                             14418 when "00110110001100",
                             14413 when "00110110001101",
                             14409 when "00110110001110",
                             14405 when "00110110001111",
                             14401 when "00110110010000",
                             14397 when "00110110010001",
                             14393 when "00110110010010",
                             14388 when "00110110010011",
                             14384 when "00110110010100",
                             14380 when "00110110010101",
                             14376 when "00110110010110",
                             14372 when "00110110010111",
                             14368 when "00110110011000",
                             14364 when "00110110011001",
                             14360 when "00110110011010",
                             14355 when "00110110011011",
                             14351 when "00110110011100",
                             14347 when "00110110011101",
                             14343 when "00110110011110",
                             14339 when "00110110011111",
                             14335 when "00110110100000",
                             14331 when "00110110100001",
                             14327 when "00110110100010",
                             14323 when "00110110100011",
                             14318 when "00110110100100",
                             14314 when "00110110100101",
                             14310 when "00110110100110",
                             14306 when "00110110100111",
                             14302 when "00110110101000",
                             14298 when "00110110101001",
                             14294 when "00110110101010",
                             14290 when "00110110101011",
                             14286 when "00110110101100",
                             14282 when "00110110101101",
                             14278 when "00110110101110",
                             14273 when "00110110101111",
                             14269 when "00110110110000",
                             14265 when "00110110110001",
                             14261 when "00110110110010",
                             14257 when "00110110110011",
                             14253 when "00110110110100",
                             14249 when "00110110110101",
                             14245 when "00110110110110",
                             14241 when "00110110110111",
                             14237 when "00110110111000",
                             14233 when "00110110111001",
                             14229 when "00110110111010",
                             14225 when "00110110111011",
                             14221 when "00110110111100",
                             14217 when "00110110111101",
                             14213 when "00110110111110",
                             14209 when "00110110111111",
                             14205 when "00110111000000",
                             14201 when "00110111000001",
                             14196 when "00110111000010",
                             14192 when "00110111000011",
                             14188 when "00110111000100",
                             14184 when "00110111000101",
                             14180 when "00110111000110",
                             14176 when "00110111000111",
                             14172 when "00110111001000",
                             14168 when "00110111001001",
                             14164 when "00110111001010",
                             14160 when "00110111001011",
                             14156 when "00110111001100",
                             14152 when "00110111001101",
                             14148 when "00110111001110",
                             14144 when "00110111001111",
                             14140 when "00110111010000",
                             14136 when "00110111010001",
                             14132 when "00110111010010",
                             14128 when "00110111010011",
                             14124 when "00110111010100",
                             14120 when "00110111010101",
                             14116 when "00110111010110",
                             14112 when "00110111010111",
                             14108 when "00110111011000",
                             14104 when "00110111011001",
                             14100 when "00110111011010",
                             14096 when "00110111011011",
                             14092 when "00110111011100",
                             14088 when "00110111011101",
                             14085 when "00110111011110",
                             14081 when "00110111011111",
                             14077 when "00110111100000",
                             14073 when "00110111100001",
                             14069 when "00110111100010",
                             14065 when "00110111100011",
                             14061 when "00110111100100",
                             14057 when "00110111100101",
                             14053 when "00110111100110",
                             14049 when "00110111100111",
                             14045 when "00110111101000",
                             14041 when "00110111101001",
                             14037 when "00110111101010",
                             14033 when "00110111101011",
                             14029 when "00110111101100",
                             14025 when "00110111101101",
                             14021 when "00110111101110",
                             14017 when "00110111101111",
                             14013 when "00110111110000",
                             14010 when "00110111110001",
                             14006 when "00110111110010",
                             14002 when "00110111110011",
                             13998 when "00110111110100",
                             13994 when "00110111110101",
                             13990 when "00110111110110",
                             13986 when "00110111110111",
                             13982 when "00110111111000",
                             13978 when "00110111111001",
                             13974 when "00110111111010",
                             13970 when "00110111111011",
                             13966 when "00110111111100",
                             13963 when "00110111111101",
                             13959 when "00110111111110",
                             13955 when "00110111111111",
                             13951 when "00111000000000",
                             13947 when "00111000000001",
                             13943 when "00111000000010",
                             13939 when "00111000000011",
                             13935 when "00111000000100",
                             13931 when "00111000000101",
                             13928 when "00111000000110",
                             13924 when "00111000000111",
                             13920 when "00111000001000",
                             13916 when "00111000001001",
                             13912 when "00111000001010",
                             13908 when "00111000001011",
                             13904 when "00111000001100",
                             13900 when "00111000001101",
                             13897 when "00111000001110",
                             13893 when "00111000001111",
                             13889 when "00111000010000",
                             13885 when "00111000010001",
                             13881 when "00111000010010",
                             13877 when "00111000010011",
                             13873 when "00111000010100",
                             13870 when "00111000010101",
                             13866 when "00111000010110",
                             13862 when "00111000010111",
                             13858 when "00111000011000",
                             13854 when "00111000011001",
                             13850 when "00111000011010",
                             13847 when "00111000011011",
                             13843 when "00111000011100",
                             13839 when "00111000011101",
                             13835 when "00111000011110",
                             13831 when "00111000011111",
                             13827 when "00111000100000",
                             13824 when "00111000100001",
                             13820 when "00111000100010",
                             13816 when "00111000100011",
                             13812 when "00111000100100",
                             13808 when "00111000100101",
                             13805 when "00111000100110",
                             13801 when "00111000100111",
                             13797 when "00111000101000",
                             13793 when "00111000101001",
                             13789 when "00111000101010",
                             13785 when "00111000101011",
                             13782 when "00111000101100",
                             13778 when "00111000101101",
                             13774 when "00111000101110",
                             13770 when "00111000101111",
                             13767 when "00111000110000",
                             13763 when "00111000110001",
                             13759 when "00111000110010",
                             13755 when "00111000110011",
                             13751 when "00111000110100",
                             13748 when "00111000110101",
                             13744 when "00111000110110",
                             13740 when "00111000110111",
                             13736 when "00111000111000",
                             13732 when "00111000111001",
                             13729 when "00111000111010",
                             13725 when "00111000111011",
                             13721 when "00111000111100",
                             13717 when "00111000111101",
                             13714 when "00111000111110",
                             13710 when "00111000111111",
                             13706 when "00111001000000",
                             13702 when "00111001000001",
                             13699 when "00111001000010",
                             13695 when "00111001000011",
                             13691 when "00111001000100",
                             13687 when "00111001000101",
                             13684 when "00111001000110",
                             13680 when "00111001000111",
                             13676 when "00111001001000",
                             13672 when "00111001001001",
                             13669 when "00111001001010",
                             13665 when "00111001001011",
                             13661 when "00111001001100",
                             13657 when "00111001001101",
                             13654 when "00111001001110",
                             13650 when "00111001001111",
                             13646 when "00111001010000",
                             13643 when "00111001010001",
                             13639 when "00111001010010",
                             13635 when "00111001010011",
                             13631 when "00111001010100",
                             13628 when "00111001010101",
                             13624 when "00111001010110",
                             13620 when "00111001010111",
                             13617 when "00111001011000",
                             13613 when "00111001011001",
                             13609 when "00111001011010",
                             13605 when "00111001011011",
                             13602 when "00111001011100",
                             13598 when "00111001011101",
                             13594 when "00111001011110",
                             13591 when "00111001011111",
                             13587 when "00111001100000",
                             13583 when "00111001100001",
                             13580 when "00111001100010",
                             13576 when "00111001100011",
                             13572 when "00111001100100",
                             13569 when "00111001100101",
                             13565 when "00111001100110",
                             13561 when "00111001100111",
                             13557 when "00111001101000",
                             13554 when "00111001101001",
                             13550 when "00111001101010",
                             13546 when "00111001101011",
                             13543 when "00111001101100",
                             13539 when "00111001101101",
                             13535 when "00111001101110",
                             13532 when "00111001101111",
                             13528 when "00111001110000",
                             13524 when "00111001110001",
                             13521 when "00111001110010",
                             13517 when "00111001110011",
                             13514 when "00111001110100",
                             13510 when "00111001110101",
                             13506 when "00111001110110",
                             13503 when "00111001110111",
                             13499 when "00111001111000",
                             13495 when "00111001111001",
                             13492 when "00111001111010",
                             13488 when "00111001111011",
                             13484 when "00111001111100",
                             13481 when "00111001111101",
                             13477 when "00111001111110",
                             13473 when "00111001111111",
                             13470 when "00111010000000",
                             13466 when "00111010000001",
                             13463 when "00111010000010",
                             13459 when "00111010000011",
                             13455 when "00111010000100",
                             13452 when "00111010000101",
                             13448 when "00111010000110",
                             13444 when "00111010000111",
                             13441 when "00111010001000",
                             13437 when "00111010001001",
                             13434 when "00111010001010",
                             13430 when "00111010001011",
                             13426 when "00111010001100",
                             13423 when "00111010001101",
                             13419 when "00111010001110",
                             13416 when "00111010001111",
                             13412 when "00111010010000",
                             13408 when "00111010010001",
                             13405 when "00111010010010",
                             13401 when "00111010010011",
                             13398 when "00111010010100",
                             13394 when "00111010010101",
                             13390 when "00111010010110",
                             13387 when "00111010010111",
                             13383 when "00111010011000",
                             13380 when "00111010011001",
                             13376 when "00111010011010",
                             13373 when "00111010011011",
                             13369 when "00111010011100",
                             13365 when "00111010011101",
                             13362 when "00111010011110",
                             13358 when "00111010011111",
                             13355 when "00111010100000",
                             13351 when "00111010100001",
                             13348 when "00111010100010",
                             13344 when "00111010100011",
                             13340 when "00111010100100",
                             13337 when "00111010100101",
                             13333 when "00111010100110",
                             13330 when "00111010100111",
                             13326 when "00111010101000",
                             13323 when "00111010101001",
                             13319 when "00111010101010",
                             13316 when "00111010101011",
                             13312 when "00111010101100",
                             13308 when "00111010101101",
                             13305 when "00111010101110",
                             13301 when "00111010101111",
                             13298 when "00111010110000",
                             13294 when "00111010110001",
                             13291 when "00111010110010",
                             13287 when "00111010110011",
                             13284 when "00111010110100",
                             13280 when "00111010110101",
                             13277 when "00111010110110",
                             13273 when "00111010110111",
                             13270 when "00111010111000",
                             13266 when "00111010111001",
                             13263 when "00111010111010",
                             13259 when "00111010111011",
                             13256 when "00111010111100",
                             13252 when "00111010111101",
                             13249 when "00111010111110",
                             13245 when "00111010111111",
                             13242 when "00111011000000",
                             13238 when "00111011000001",
                             13235 when "00111011000010",
                             13231 when "00111011000011",
                             13228 when "00111011000100",
                             13224 when "00111011000101",
                             13221 when "00111011000110",
                             13217 when "00111011000111",
                             13214 when "00111011001000",
                             13210 when "00111011001001",
                             13207 when "00111011001010",
                             13203 when "00111011001011",
                             13200 when "00111011001100",
                             13196 when "00111011001101",
                             13193 when "00111011001110",
                             13189 when "00111011001111",
                             13186 when "00111011010000",
                             13182 when "00111011010001",
                             13179 when "00111011010010",
                             13175 when "00111011010011",
                             13172 when "00111011010100",
                             13168 when "00111011010101",
                             13165 when "00111011010110",
                             13161 when "00111011010111",
                             13158 when "00111011011000",
                             13154 when "00111011011001",
                             13151 when "00111011011010",
                             13148 when "00111011011011",
                             13144 when "00111011011100",
                             13141 when "00111011011101",
                             13137 when "00111011011110",
                             13134 when "00111011011111",
                             13130 when "00111011100000",
                             13127 when "00111011100001",
                             13123 when "00111011100010",
                             13120 when "00111011100011",
                             13116 when "00111011100100",
                             13113 when "00111011100101",
                             13110 when "00111011100110",
                             13106 when "00111011100111",
                             13103 when "00111011101000",
                             13099 when "00111011101001",
                             13096 when "00111011101010",
                             13092 when "00111011101011",
                             13089 when "00111011101100",
                             13086 when "00111011101101",
                             13082 when "00111011101110",
                             13079 when "00111011101111",
                             13075 when "00111011110000",
                             13072 when "00111011110001",
                             13068 when "00111011110010",
                             13065 when "00111011110011",
                             13062 when "00111011110100",
                             13058 when "00111011110101",
                             13055 when "00111011110110",
                             13051 when "00111011110111",
                             13048 when "00111011111000",
                             13045 when "00111011111001",
                             13041 when "00111011111010",
                             13038 when "00111011111011",
                             13034 when "00111011111100",
                             13031 when "00111011111101",
                             13028 when "00111011111110",
                             13024 when "00111011111111",
                             13021 when "00111100000000",
                             13017 when "00111100000001",
                             13014 when "00111100000010",
                             13011 when "00111100000011",
                             13007 when "00111100000100",
                             13004 when "00111100000101",
                             13001 when "00111100000110",
                             12997 when "00111100000111",
                             12994 when "00111100001000",
                             12990 when "00111100001001",
                             12987 when "00111100001010",
                             12984 when "00111100001011",
                             12980 when "00111100001100",
                             12977 when "00111100001101",
                             12974 when "00111100001110",
                             12970 when "00111100001111",
                             12967 when "00111100010000",
                             12963 when "00111100010001",
                             12960 when "00111100010010",
                             12957 when "00111100010011",
                             12953 when "00111100010100",
                             12950 when "00111100010101",
                             12947 when "00111100010110",
                             12943 when "00111100010111",
                             12940 when "00111100011000",
                             12937 when "00111100011001",
                             12933 when "00111100011010",
                             12930 when "00111100011011",
                             12927 when "00111100011100",
                             12923 when "00111100011101",
                             12920 when "00111100011110",
                             12917 when "00111100011111",
                             12913 when "00111100100000",
                             12910 when "00111100100001",
                             12907 when "00111100100010",
                             12903 when "00111100100011",
                             12900 when "00111100100100",
                             12897 when "00111100100101",
                             12893 when "00111100100110",
                             12890 when "00111100100111",
                             12887 when "00111100101000",
                             12883 when "00111100101001",
                             12880 when "00111100101010",
                             12877 when "00111100101011",
                             12873 when "00111100101100",
                             12870 when "00111100101101",
                             12867 when "00111100101110",
                             12863 when "00111100101111",
                             12860 when "00111100110000",
                             12857 when "00111100110001",
                             12853 when "00111100110010",
                             12850 when "00111100110011",
                             12847 when "00111100110100",
                             12844 when "00111100110101",
                             12840 when "00111100110110",
                             12837 when "00111100110111",
                             12834 when "00111100111000",
                             12830 when "00111100111001",
                             12827 when "00111100111010",
                             12824 when "00111100111011",
                             12821 when "00111100111100",
                             12817 when "00111100111101",
                             12814 when "00111100111110",
                             12811 when "00111100111111",
                             12807 when "00111101000000",
                             12804 when "00111101000001",
                             12801 when "00111101000010",
                             12798 when "00111101000011",
                             12794 when "00111101000100",
                             12791 when "00111101000101",
                             12788 when "00111101000110",
                             12784 when "00111101000111",
                             12781 when "00111101001000",
                             12778 when "00111101001001",
                             12775 when "00111101001010",
                             12771 when "00111101001011",
                             12768 when "00111101001100",
                             12765 when "00111101001101",
                             12762 when "00111101001110",
                             12758 when "00111101001111",
                             12755 when "00111101010000",
                             12752 when "00111101010001",
                             12749 when "00111101010010",
                             12745 when "00111101010011",
                             12742 when "00111101010100",
                             12739 when "00111101010101",
                             12736 when "00111101010110",
                             12732 when "00111101010111",
                             12729 when "00111101011000",
                             12726 when "00111101011001",
                             12723 when "00111101011010",
                             12719 when "00111101011011",
                             12716 when "00111101011100",
                             12713 when "00111101011101",
                             12710 when "00111101011110",
                             12706 when "00111101011111",
                             12703 when "00111101100000",
                             12700 when "00111101100001",
                             12697 when "00111101100010",
                             12694 when "00111101100011",
                             12690 when "00111101100100",
                             12687 when "00111101100101",
                             12684 when "00111101100110",
                             12681 when "00111101100111",
                             12677 when "00111101101000",
                             12674 when "00111101101001",
                             12671 when "00111101101010",
                             12668 when "00111101101011",
                             12665 when "00111101101100",
                             12661 when "00111101101101",
                             12658 when "00111101101110",
                             12655 when "00111101101111",
                             12652 when "00111101110000",
                             12649 when "00111101110001",
                             12645 when "00111101110010",
                             12642 when "00111101110011",
                             12639 when "00111101110100",
                             12636 when "00111101110101",
                             12633 when "00111101110110",
                             12629 when "00111101110111",
                             12626 when "00111101111000",
                             12623 when "00111101111001",
                             12620 when "00111101111010",
                             12617 when "00111101111011",
                             12614 when "00111101111100",
                             12610 when "00111101111101",
                             12607 when "00111101111110",
                             12604 when "00111101111111",
                             12601 when "00111110000000",
                             12598 when "00111110000001",
                             12594 when "00111110000010",
                             12591 when "00111110000011",
                             12588 when "00111110000100",
                             12585 when "00111110000101",
                             12582 when "00111110000110",
                             12579 when "00111110000111",
                             12575 when "00111110001000",
                             12572 when "00111110001001",
                             12569 when "00111110001010",
                             12566 when "00111110001011",
                             12563 when "00111110001100",
                             12560 when "00111110001101",
                             12557 when "00111110001110",
                             12553 when "00111110001111",
                             12550 when "00111110010000",
                             12547 when "00111110010001",
                             12544 when "00111110010010",
                             12541 when "00111110010011",
                             12538 when "00111110010100",
                             12534 when "00111110010101",
                             12531 when "00111110010110",
                             12528 when "00111110010111",
                             12525 when "00111110011000",
                             12522 when "00111110011001",
                             12519 when "00111110011010",
                             12516 when "00111110011011",
                             12513 when "00111110011100",
                             12509 when "00111110011101",
                             12506 when "00111110011110",
                             12503 when "00111110011111",
                             12500 when "00111110100000",
                             12497 when "00111110100001",
                             12494 when "00111110100010",
                             12491 when "00111110100011",
                             12488 when "00111110100100",
                             12484 when "00111110100101",
                             12481 when "00111110100110",
                             12478 when "00111110100111",
                             12475 when "00111110101000",
                             12472 when "00111110101001",
                             12469 when "00111110101010",
                             12466 when "00111110101011",
                             12463 when "00111110101100",
                             12460 when "00111110101101",
                             12456 when "00111110101110",
                             12453 when "00111110101111",
                             12450 when "00111110110000",
                             12447 when "00111110110001",
                             12444 when "00111110110010",
                             12441 when "00111110110011",
                             12438 when "00111110110100",
                             12435 when "00111110110101",
                             12432 when "00111110110110",
                             12429 when "00111110110111",
                             12425 when "00111110111000",
                             12422 when "00111110111001",
                             12419 when "00111110111010",
                             12416 when "00111110111011",
                             12413 when "00111110111100",
                             12410 when "00111110111101",
                             12407 when "00111110111110",
                             12404 when "00111110111111",
                             12401 when "00111111000000",
                             12398 when "00111111000001",
                             12395 when "00111111000010",
                             12392 when "00111111000011",
                             12389 when "00111111000100",
                             12385 when "00111111000101",
                             12382 when "00111111000110",
                             12379 when "00111111000111",
                             12376 when "00111111001000",
                             12373 when "00111111001001",
                             12370 when "00111111001010",
                             12367 when "00111111001011",
                             12364 when "00111111001100",
                             12361 when "00111111001101",
                             12358 when "00111111001110",
                             12355 when "00111111001111",
                             12352 when "00111111010000",
                             12349 when "00111111010001",
                             12346 when "00111111010010",
                             12343 when "00111111010011",
                             12340 when "00111111010100",
                             12337 when "00111111010101",
                             12333 when "00111111010110",
                             12330 when "00111111010111",
                             12327 when "00111111011000",
                             12324 when "00111111011001",
                             12321 when "00111111011010",
                             12318 when "00111111011011",
                             12315 when "00111111011100",
                             12312 when "00111111011101",
                             12309 when "00111111011110",
                             12306 when "00111111011111",
                             12303 when "00111111100000",
                             12300 when "00111111100001",
                             12297 when "00111111100010",
                             12294 when "00111111100011",
                             12291 when "00111111100100",
                             12288 when "00111111100101",
                             12285 when "00111111100110",
                             12282 when "00111111100111",
                             12279 when "00111111101000",
                             12276 when "00111111101001",
                             12273 when "00111111101010",
                             12270 when "00111111101011",
                             12267 when "00111111101100",
                             12264 when "00111111101101",
                             12261 when "00111111101110",
                             12258 when "00111111101111",
                             12255 when "00111111110000",
                             12252 when "00111111110001",
                             12249 when "00111111110010",
                             12246 when "00111111110011",
                             12243 when "00111111110100",
                             12240 when "00111111110101",
                             12237 when "00111111110110",
                             12234 when "00111111110111",
                             12231 when "00111111111000",
                             12228 when "00111111111001",
                             12225 when "00111111111010",
                             12222 when "00111111111011",
                             12219 when "00111111111100",
                             12216 when "00111111111101",
                             12213 when "00111111111110",
                             12210 when "00111111111111",
                             12207 when "01000000000000",
                             12204 when "01000000000001",
                             12201 when "01000000000010",
                             12198 when "01000000000011",
                             12195 when "01000000000100",
                             12192 when "01000000000101",
                             12189 when "01000000000110",
                             12186 when "01000000000111",
                             12183 when "01000000001000",
                             12180 when "01000000001001",
                             12177 when "01000000001010",
                             12174 when "01000000001011",
                             12171 when "01000000001100",
                             12168 when "01000000001101",
                             12165 when "01000000001110",
                             12162 when "01000000001111",
                             12160 when "01000000010000",
                             12157 when "01000000010001",
                             12154 when "01000000010010",
                             12151 when "01000000010011",
                             12148 when "01000000010100",
                             12145 when "01000000010101",
                             12142 when "01000000010110",
                             12139 when "01000000010111",
                             12136 when "01000000011000",
                             12133 when "01000000011001",
                             12130 when "01000000011010",
                             12127 when "01000000011011",
                             12124 when "01000000011100",
                             12121 when "01000000011101",
                             12118 when "01000000011110",
                             12115 when "01000000011111",
                             12112 when "01000000100000",
                             12109 when "01000000100001",
                             12107 when "01000000100010",
                             12104 when "01000000100011",
                             12101 when "01000000100100",
                             12098 when "01000000100101",
                             12095 when "01000000100110",
                             12092 when "01000000100111",
                             12089 when "01000000101000",
                             12086 when "01000000101001",
                             12083 when "01000000101010",
                             12080 when "01000000101011",
                             12077 when "01000000101100",
                             12074 when "01000000101101",
                             12071 when "01000000101110",
                             12069 when "01000000101111",
                             12066 when "01000000110000",
                             12063 when "01000000110001",
                             12060 when "01000000110010",
                             12057 when "01000000110011",
                             12054 when "01000000110100",
                             12051 when "01000000110101",
                             12048 when "01000000110110",
                             12045 when "01000000110111",
                             12042 when "01000000111000",
                             12039 when "01000000111001",
                             12037 when "01000000111010",
                             12034 when "01000000111011",
                             12031 when "01000000111100",
                             12028 when "01000000111101",
                             12025 when "01000000111110",
                             12022 when "01000000111111",
                             12019 when "01000001000000",
                             12016 when "01000001000001",
                             12013 when "01000001000010",
                             12011 when "01000001000011",
                             12008 when "01000001000100",
                             12005 when "01000001000101",
                             12002 when "01000001000110",
                             11999 when "01000001000111",
                             11996 when "01000001001000",
                             11993 when "01000001001001",
                             11990 when "01000001001010",
                             11988 when "01000001001011",
                             11985 when "01000001001100",
                             11982 when "01000001001101",
                             11979 when "01000001001110",
                             11976 when "01000001001111",
                             11973 when "01000001010000",
                             11970 when "01000001010001",
                             11967 when "01000001010010",
                             11965 when "01000001010011",
                             11962 when "01000001010100",
                             11959 when "01000001010101",
                             11956 when "01000001010110",
                             11953 when "01000001010111",
                             11950 when "01000001011000",
                             11947 when "01000001011001",
                             11945 when "01000001011010",
                             11942 when "01000001011011",
                             11939 when "01000001011100",
                             11936 when "01000001011101",
                             11933 when "01000001011110",
                             11930 when "01000001011111",
                             11927 when "01000001100000",
                             11925 when "01000001100001",
                             11922 when "01000001100010",
                             11919 when "01000001100011",
                             11916 when "01000001100100",
                             11913 when "01000001100101",
                             11910 when "01000001100110",
                             11908 when "01000001100111",
                             11905 when "01000001101000",
                             11902 when "01000001101001",
                             11899 when "01000001101010",
                             11896 when "01000001101011",
                             11893 when "01000001101100",
                             11891 when "01000001101101",
                             11888 when "01000001101110",
                             11885 when "01000001101111",
                             11882 when "01000001110000",
                             11879 when "01000001110001",
                             11876 when "01000001110010",
                             11874 when "01000001110011",
                             11871 when "01000001110100",
                             11868 when "01000001110101",
                             11865 when "01000001110110",
                             11862 when "01000001110111",
                             11860 when "01000001111000",
                             11857 when "01000001111001",
                             11854 when "01000001111010",
                             11851 when "01000001111011",
                             11848 when "01000001111100",
                             11846 when "01000001111101",
                             11843 when "01000001111110",
                             11840 when "01000001111111",
                             11837 when "01000010000000",
                             11834 when "01000010000001",
                             11832 when "01000010000010",
                             11829 when "01000010000011",
                             11826 when "01000010000100",
                             11823 when "01000010000101",
                             11820 when "01000010000110",
                             11818 when "01000010000111",
                             11815 when "01000010001000",
                             11812 when "01000010001001",
                             11809 when "01000010001010",
                             11806 when "01000010001011",
                             11804 when "01000010001100",
                             11801 when "01000010001101",
                             11798 when "01000010001110",
                             11795 when "01000010001111",
                             11792 when "01000010010000",
                             11790 when "01000010010001",
                             11787 when "01000010010010",
                             11784 when "01000010010011",
                             11781 when "01000010010100",
                             11779 when "01000010010101",
                             11776 when "01000010010110",
                             11773 when "01000010010111",
                             11770 when "01000010011000",
                             11767 when "01000010011001",
                             11765 when "01000010011010",
                             11762 when "01000010011011",
                             11759 when "01000010011100",
                             11756 when "01000010011101",
                             11754 when "01000010011110",
                             11751 when "01000010011111",
                             11748 when "01000010100000",
                             11745 when "01000010100001",
                             11743 when "01000010100010",
                             11740 when "01000010100011",
                             11737 when "01000010100100",
                             11734 when "01000010100101",
                             11732 when "01000010100110",
                             11729 when "01000010100111",
                             11726 when "01000010101000",
                             11723 when "01000010101001",
                             11721 when "01000010101010",
                             11718 when "01000010101011",
                             11715 when "01000010101100",
                             11712 when "01000010101101",
                             11710 when "01000010101110",
                             11707 when "01000010101111",
                             11704 when "01000010110000",
                             11701 when "01000010110001",
                             11699 when "01000010110010",
                             11696 when "01000010110011",
                             11693 when "01000010110100",
                             11690 when "01000010110101",
                             11688 when "01000010110110",
                             11685 when "01000010110111",
                             11682 when "01000010111000",
                             11680 when "01000010111001",
                             11677 when "01000010111010",
                             11674 when "01000010111011",
                             11671 when "01000010111100",
                             11669 when "01000010111101",
                             11666 when "01000010111110",
                             11663 when "01000010111111",
                             11660 when "01000011000000",
                             11658 when "01000011000001",
                             11655 when "01000011000010",
                             11652 when "01000011000011",
                             11650 when "01000011000100",
                             11647 when "01000011000101",
                             11644 when "01000011000110",
                             11641 when "01000011000111",
                             11639 when "01000011001000",
                             11636 when "01000011001001",
                             11633 when "01000011001010",
                             11631 when "01000011001011",
                             11628 when "01000011001100",
                             11625 when "01000011001101",
                             11623 when "01000011001110",
                             11620 when "01000011001111",
                             11617 when "01000011010000",
                             11614 when "01000011010001",
                             11612 when "01000011010010",
                             11609 when "01000011010011",
                             11606 when "01000011010100",
                             11604 when "01000011010101",
                             11601 when "01000011010110",
                             11598 when "01000011010111",
                             11596 when "01000011011000",
                             11593 when "01000011011001",
                             11590 when "01000011011010",
                             11587 when "01000011011011",
                             11585 when "01000011011100",
                             11582 when "01000011011101",
                             11579 when "01000011011110",
                             11577 when "01000011011111",
                             11574 when "01000011100000",
                             11571 when "01000011100001",
                             11569 when "01000011100010",
                             11566 when "01000011100011",
                             11563 when "01000011100100",
                             11561 when "01000011100101",
                             11558 when "01000011100110",
                             11555 when "01000011100111",
                             11553 when "01000011101000",
                             11550 when "01000011101001",
                             11547 when "01000011101010",
                             11545 when "01000011101011",
                             11542 when "01000011101100",
                             11539 when "01000011101101",
                             11537 when "01000011101110",
                             11534 when "01000011101111",
                             11531 when "01000011110000",
                             11529 when "01000011110001",
                             11526 when "01000011110010",
                             11523 when "01000011110011",
                             11521 when "01000011110100",
                             11518 when "01000011110101",
                             11515 when "01000011110110",
                             11513 when "01000011110111",
                             11510 when "01000011111000",
                             11507 when "01000011111001",
                             11505 when "01000011111010",
                             11502 when "01000011111011",
                             11500 when "01000011111100",
                             11497 when "01000011111101",
                             11494 when "01000011111110",
                             11492 when "01000011111111",
                             11489 when "01000100000000",
                             11486 when "01000100000001",
                             11484 when "01000100000010",
                             11481 when "01000100000011",
                             11478 when "01000100000100",
                             11476 when "01000100000101",
                             11473 when "01000100000110",
                             11471 when "01000100000111",
                             11468 when "01000100001000",
                             11465 when "01000100001001",
                             11463 when "01000100001010",
                             11460 when "01000100001011",
                             11457 when "01000100001100",
                             11455 when "01000100001101",
                             11452 when "01000100001110",
                             11450 when "01000100001111",
                             11447 when "01000100010000",
                             11444 when "01000100010001",
                             11442 when "01000100010010",
                             11439 when "01000100010011",
                             11436 when "01000100010100",
                             11434 when "01000100010101",
                             11431 when "01000100010110",
                             11429 when "01000100010111",
                             11426 when "01000100011000",
                             11423 when "01000100011001",
                             11421 when "01000100011010",
                             11418 when "01000100011011",
                             11416 when "01000100011100",
                             11413 when "01000100011101",
                             11410 when "01000100011110",
                             11408 when "01000100011111",
                             11405 when "01000100100000",
                             11403 when "01000100100001",
                             11400 when "01000100100010",
                             11397 when "01000100100011",
                             11395 when "01000100100100",
                             11392 when "01000100100101",
                             11390 when "01000100100110",
                             11387 when "01000100100111",
                             11384 when "01000100101000",
                             11382 when "01000100101001",
                             11379 when "01000100101010",
                             11377 when "01000100101011",
                             11374 when "01000100101100",
                             11371 when "01000100101101",
                             11369 when "01000100101110",
                             11366 when "01000100101111",
                             11364 when "01000100110000",
                             11361 when "01000100110001",
                             11358 when "01000100110010",
                             11356 when "01000100110011",
                             11353 when "01000100110100",
                             11351 when "01000100110101",
                             11348 when "01000100110110",
                             11346 when "01000100110111",
                             11343 when "01000100111000",
                             11340 when "01000100111001",
                             11338 when "01000100111010",
                             11335 when "01000100111011",
                             11333 when "01000100111100",
                             11330 when "01000100111101",
                             11328 when "01000100111110",
                             11325 when "01000100111111",
                             11322 when "01000101000000",
                             11320 when "01000101000001",
                             11317 when "01000101000010",
                             11315 when "01000101000011",
                             11312 when "01000101000100",
                             11310 when "01000101000101",
                             11307 when "01000101000110",
                             11305 when "01000101000111",
                             11302 when "01000101001000",
                             11299 when "01000101001001",
                             11297 when "01000101001010",
                             11294 when "01000101001011",
                             11292 when "01000101001100",
                             11289 when "01000101001101",
                             11287 when "01000101001110",
                             11284 when "01000101001111",
                             11282 when "01000101010000",
                             11279 when "01000101010001",
                             11276 when "01000101010010",
                             11274 when "01000101010011",
                             11271 when "01000101010100",
                             11269 when "01000101010101",
                             11266 when "01000101010110",
                             11264 when "01000101010111",
                             11261 when "01000101011000",
                             11259 when "01000101011001",
                             11256 when "01000101011010",
                             11254 when "01000101011011",
                             11251 when "01000101011100",
                             11249 when "01000101011101",
                             11246 when "01000101011110",
                             11244 when "01000101011111",
                             11241 when "01000101100000",
                             11238 when "01000101100001",
                             11236 when "01000101100010",
                             11233 when "01000101100011",
                             11231 when "01000101100100",
                             11228 when "01000101100101",
                             11226 when "01000101100110",
                             11223 when "01000101100111",
                             11221 when "01000101101000",
                             11218 when "01000101101001",
                             11216 when "01000101101010",
                             11213 when "01000101101011",
                             11211 when "01000101101100",
                             11208 when "01000101101101",
                             11206 when "01000101101110",
                             11203 when "01000101101111",
                             11201 when "01000101110000",
                             11198 when "01000101110001",
                             11196 when "01000101110010",
                             11193 when "01000101110011",
                             11191 when "01000101110100",
                             11188 when "01000101110101",
                             11186 when "01000101110110",
                             11183 when "01000101110111",
                             11181 when "01000101111000",
                             11178 when "01000101111001",
                             11176 when "01000101111010",
                             11173 when "01000101111011",
                             11171 when "01000101111100",
                             11168 when "01000101111101",
                             11166 when "01000101111110",
                             11163 when "01000101111111",
                             11161 when "01000110000000",
                             11158 when "01000110000001",
                             11156 when "01000110000010",
                             11153 when "01000110000011",
                             11151 when "01000110000100",
                             11148 when "01000110000101",
                             11146 when "01000110000110",
                             11143 when "01000110000111",
                             11141 when "01000110001000",
                             11138 when "01000110001001",
                             11136 when "01000110001010",
                             11133 when "01000110001011",
                             11131 when "01000110001100",
                             11128 when "01000110001101",
                             11126 when "01000110001110",
                             11123 when "01000110001111",
                             11121 when "01000110010000",
                             11119 when "01000110010001",
                             11116 when "01000110010010",
                             11114 when "01000110010011",
                             11111 when "01000110010100",
                             11109 when "01000110010101",
                             11106 when "01000110010110",
                             11104 when "01000110010111",
                             11101 when "01000110011000",
                             11099 when "01000110011001",
                             11096 when "01000110011010",
                             11094 when "01000110011011",
                             11091 when "01000110011100",
                             11089 when "01000110011101",
                             11086 when "01000110011110",
                             11084 when "01000110011111",
                             11082 when "01000110100000",
                             11079 when "01000110100001",
                             11077 when "01000110100010",
                             11074 when "01000110100011",
                             11072 when "01000110100100",
                             11069 when "01000110100101",
                             11067 when "01000110100110",
                             11064 when "01000110100111",
                             11062 when "01000110101000",
                             11060 when "01000110101001",
                             11057 when "01000110101010",
                             11055 when "01000110101011",
                             11052 when "01000110101100",
                             11050 when "01000110101101",
                             11047 when "01000110101110",
                             11045 when "01000110101111",
                             11042 when "01000110110000",
                             11040 when "01000110110001",
                             11038 when "01000110110010",
                             11035 when "01000110110011",
                             11033 when "01000110110100",
                             11030 when "01000110110101",
                             11028 when "01000110110110",
                             11025 when "01000110110111",
                             11023 when "01000110111000",
                             11020 when "01000110111001",
                             11018 when "01000110111010",
                             11016 when "01000110111011",
                             11013 when "01000110111100",
                             11011 when "01000110111101",
                             11008 when "01000110111110",
                             11006 when "01000110111111",
                             11004 when "01000111000000",
                             11001 when "01000111000001",
                             10999 when "01000111000010",
                             10996 when "01000111000011",
                             10994 when "01000111000100",
                             10991 when "01000111000101",
                             10989 when "01000111000110",
                             10987 when "01000111000111",
                             10984 when "01000111001000",
                             10982 when "01000111001001",
                             10979 when "01000111001010",
                             10977 when "01000111001011",
                             10975 when "01000111001100",
                             10972 when "01000111001101",
                             10970 when "01000111001110",
                             10967 when "01000111001111",
                             10965 when "01000111010000",
                             10963 when "01000111010001",
                             10960 when "01000111010010",
                             10958 when "01000111010011",
                             10955 when "01000111010100",
                             10953 when "01000111010101",
                             10951 when "01000111010110",
                             10948 when "01000111010111",
                             10946 when "01000111011000",
                             10943 when "01000111011001",
                             10941 when "01000111011010",
                             10939 when "01000111011011",
                             10936 when "01000111011100",
                             10934 when "01000111011101",
                             10931 when "01000111011110",
                             10929 when "01000111011111",
                             10927 when "01000111100000",
                             10924 when "01000111100001",
                             10922 when "01000111100010",
                             10919 when "01000111100011",
                             10917 when "01000111100100",
                             10915 when "01000111100101",
                             10912 when "01000111100110",
                             10910 when "01000111100111",
                             10908 when "01000111101000",
                             10905 when "01000111101001",
                             10903 when "01000111101010",
                             10900 when "01000111101011",
                             10898 when "01000111101100",
                             10896 when "01000111101101",
                             10893 when "01000111101110",
                             10891 when "01000111101111",
                             10889 when "01000111110000",
                             10886 when "01000111110001",
                             10884 when "01000111110010",
                             10881 when "01000111110011",
                             10879 when "01000111110100",
                             10877 when "01000111110101",
                             10874 when "01000111110110",
                             10872 when "01000111110111",
                             10870 when "01000111111000",
                             10867 when "01000111111001",
                             10865 when "01000111111010",
                             10862 when "01000111111011",
                             10860 when "01000111111100",
                             10858 when "01000111111101",
                             10855 when "01000111111110",
                             10853 when "01000111111111",
                             10851 when "01001000000000",
                             10848 when "01001000000001",
                             10846 when "01001000000010",
                             10844 when "01001000000011",
                             10841 when "01001000000100",
                             10839 when "01001000000101",
                             10837 when "01001000000110",
                             10834 when "01001000000111",
                             10832 when "01001000001000",
                             10830 when "01001000001001",
                             10827 when "01001000001010",
                             10825 when "01001000001011",
                             10823 when "01001000001100",
                             10820 when "01001000001101",
                             10818 when "01001000001110",
                             10815 when "01001000001111",
                             10813 when "01001000010000",
                             10811 when "01001000010001",
                             10808 when "01001000010010",
                             10806 when "01001000010011",
                             10804 when "01001000010100",
                             10801 when "01001000010101",
                             10799 when "01001000010110",
                             10797 when "01001000010111",
                             10794 when "01001000011000",
                             10792 when "01001000011001",
                             10790 when "01001000011010",
                             10787 when "01001000011011",
                             10785 when "01001000011100",
                             10783 when "01001000011101",
                             10781 when "01001000011110",
                             10778 when "01001000011111",
                             10776 when "01001000100000",
                             10774 when "01001000100001",
                             10771 when "01001000100010",
                             10769 when "01001000100011",
                             10767 when "01001000100100",
                             10764 when "01001000100101",
                             10762 when "01001000100110",
                             10760 when "01001000100111",
                             10757 when "01001000101000",
                             10755 when "01001000101001",
                             10753 when "01001000101010",
                             10750 when "01001000101011",
                             10748 when "01001000101100",
                             10746 when "01001000101101",
                             10743 when "01001000101110",
                             10741 when "01001000101111",
                             10739 when "01001000110000",
                             10737 when "01001000110001",
                             10734 when "01001000110010",
                             10732 when "01001000110011",
                             10730 when "01001000110100",
                             10727 when "01001000110101",
                             10725 when "01001000110110",
                             10723 when "01001000110111",
                             10720 when "01001000111000",
                             10718 when "01001000111001",
                             10716 when "01001000111010",
                             10714 when "01001000111011",
                             10711 when "01001000111100",
                             10709 when "01001000111101",
                             10707 when "01001000111110",
                             10704 when "01001000111111",
                             10702 when "01001001000000",
                             10700 when "01001001000001",
                             10697 when "01001001000010",
                             10695 when "01001001000011",
                             10693 when "01001001000100",
                             10691 when "01001001000101",
                             10688 when "01001001000110",
                             10686 when "01001001000111",
                             10684 when "01001001001000",
                             10681 when "01001001001001",
                             10679 when "01001001001010",
                             10677 when "01001001001011",
                             10675 when "01001001001100",
                             10672 when "01001001001101",
                             10670 when "01001001001110",
                             10668 when "01001001001111",
                             10666 when "01001001010000",
                             10663 when "01001001010001",
                             10661 when "01001001010010",
                             10659 when "01001001010011",
                             10656 when "01001001010100",
                             10654 when "01001001010101",
                             10652 when "01001001010110",
                             10650 when "01001001010111",
                             10647 when "01001001011000",
                             10645 when "01001001011001",
                             10643 when "01001001011010",
                             10641 when "01001001011011",
                             10638 when "01001001011100",
                             10636 when "01001001011101",
                             10634 when "01001001011110",
                             10632 when "01001001011111",
                             10629 when "01001001100000",
                             10627 when "01001001100001",
                             10625 when "01001001100010",
                             10622 when "01001001100011",
                             10620 when "01001001100100",
                             10618 when "01001001100101",
                             10616 when "01001001100110",
                             10613 when "01001001100111",
                             10611 when "01001001101000",
                             10609 when "01001001101001",
                             10607 when "01001001101010",
                             10604 when "01001001101011",
                             10602 when "01001001101100",
                             10600 when "01001001101101",
                             10598 when "01001001101110",
                             10595 when "01001001101111",
                             10593 when "01001001110000",
                             10591 when "01001001110001",
                             10589 when "01001001110010",
                             10586 when "01001001110011",
                             10584 when "01001001110100",
                             10582 when "01001001110101",
                             10580 when "01001001110110",
                             10578 when "01001001110111",
                             10575 when "01001001111000",
                             10573 when "01001001111001",
                             10571 when "01001001111010",
                             10569 when "01001001111011",
                             10566 when "01001001111100",
                             10564 when "01001001111101",
                             10562 when "01001001111110",
                             10560 when "01001001111111",
                             10557 when "01001010000000",
                             10555 when "01001010000001",
                             10553 when "01001010000010",
                             10551 when "01001010000011",
                             10549 when "01001010000100",
                             10546 when "01001010000101",
                             10544 when "01001010000110",
                             10542 when "01001010000111",
                             10540 when "01001010001000",
                             10537 when "01001010001001",
                             10535 when "01001010001010",
                             10533 when "01001010001011",
                             10531 when "01001010001100",
                             10529 when "01001010001101",
                             10526 when "01001010001110",
                             10524 when "01001010001111",
                             10522 when "01001010010000",
                             10520 when "01001010010001",
                             10517 when "01001010010010",
                             10515 when "01001010010011",
                             10513 when "01001010010100",
                             10511 when "01001010010101",
                             10509 when "01001010010110",
                             10506 when "01001010010111",
                             10504 when "01001010011000",
                             10502 when "01001010011001",
                             10500 when "01001010011010",
                             10498 when "01001010011011",
                             10495 when "01001010011100",
                             10493 when "01001010011101",
                             10491 when "01001010011110",
                             10489 when "01001010011111",
                             10487 when "01001010100000",
                             10484 when "01001010100001",
                             10482 when "01001010100010",
                             10480 when "01001010100011",
                             10478 when "01001010100100",
                             10476 when "01001010100101",
                             10473 when "01001010100110",
                             10471 when "01001010100111",
                             10469 when "01001010101000",
                             10467 when "01001010101001",
                             10465 when "01001010101010",
                             10462 when "01001010101011",
                             10460 when "01001010101100",
                             10458 when "01001010101101",
                             10456 when "01001010101110",
                             10454 when "01001010101111",
                             10452 when "01001010110000",
                             10449 when "01001010110001",
                             10447 when "01001010110010",
                             10445 when "01001010110011",
                             10443 when "01001010110100",
                             10441 when "01001010110101",
                             10438 when "01001010110110",
                             10436 when "01001010110111",
                             10434 when "01001010111000",
                             10432 when "01001010111001",
                             10430 when "01001010111010",
                             10428 when "01001010111011",
                             10425 when "01001010111100",
                             10423 when "01001010111101",
                             10421 when "01001010111110",
                             10419 when "01001010111111",
                             10417 when "01001011000000",
                             10414 when "01001011000001",
                             10412 when "01001011000010",
                             10410 when "01001011000011",
                             10408 when "01001011000100",
                             10406 when "01001011000101",
                             10404 when "01001011000110",
                             10401 when "01001011000111",
                             10399 when "01001011001000",
                             10397 when "01001011001001",
                             10395 when "01001011001010",
                             10393 when "01001011001011",
                             10391 when "01001011001100",
                             10389 when "01001011001101",
                             10386 when "01001011001110",
                             10384 when "01001011001111",
                             10382 when "01001011010000",
                             10380 when "01001011010001",
                             10378 when "01001011010010",
                             10376 when "01001011010011",
                             10373 when "01001011010100",
                             10371 when "01001011010101",
                             10369 when "01001011010110",
                             10367 when "01001011010111",
                             10365 when "01001011011000",
                             10363 when "01001011011001",
                             10361 when "01001011011010",
                             10358 when "01001011011011",
                             10356 when "01001011011100",
                             10354 when "01001011011101",
                             10352 when "01001011011110",
                             10350 when "01001011011111",
                             10348 when "01001011100000",
                             10346 when "01001011100001",
                             10343 when "01001011100010",
                             10341 when "01001011100011",
                             10339 when "01001011100100",
                             10337 when "01001011100101",
                             10335 when "01001011100110",
                             10333 when "01001011100111",
                             10331 when "01001011101000",
                             10328 when "01001011101001",
                             10326 when "01001011101010",
                             10324 when "01001011101011",
                             10322 when "01001011101100",
                             10320 when "01001011101101",
                             10318 when "01001011101110",
                             10316 when "01001011101111",
                             10314 when "01001011110000",
                             10311 when "01001011110001",
                             10309 when "01001011110010",
                             10307 when "01001011110011",
                             10305 when "01001011110100",
                             10303 when "01001011110101",
                             10301 when "01001011110110",
                             10299 when "01001011110111",
                             10297 when "01001011111000",
                             10294 when "01001011111001",
                             10292 when "01001011111010",
                             10290 when "01001011111011",
                             10288 when "01001011111100",
                             10286 when "01001011111101",
                             10284 when "01001011111110",
                             10282 when "01001011111111",
                             10280 when "01001100000000",
                             10277 when "01001100000001",
                             10275 when "01001100000010",
                             10273 when "01001100000011",
                             10271 when "01001100000100",
                             10269 when "01001100000101",
                             10267 when "01001100000110",
                             10265 when "01001100000111",
                             10263 when "01001100001000",
                             10261 when "01001100001001",
                             10259 when "01001100001010",
                             10256 when "01001100001011",
                             10254 when "01001100001100",
                             10252 when "01001100001101",
                             10250 when "01001100001110",
                             10248 when "01001100001111",
                             10246 when "01001100010000",
                             10244 when "01001100010001",
                             10242 when "01001100010010",
                             10240 when "01001100010011",
                             10238 when "01001100010100",
                             10235 when "01001100010101",
                             10233 when "01001100010110",
                             10231 when "01001100010111",
                             10229 when "01001100011000",
                             10227 when "01001100011001",
                             10225 when "01001100011010",
                             10223 when "01001100011011",
                             10221 when "01001100011100",
                             10219 when "01001100011101",
                             10217 when "01001100011110",
                             10215 when "01001100011111",
                             10212 when "01001100100000",
                             10210 when "01001100100001",
                             10208 when "01001100100010",
                             10206 when "01001100100011",
                             10204 when "01001100100100",
                             10202 when "01001100100101",
                             10200 when "01001100100110",
                             10198 when "01001100100111",
                             10196 when "01001100101000",
                             10194 when "01001100101001",
                             10192 when "01001100101010",
                             10190 when "01001100101011",
                             10187 when "01001100101100",
                             10185 when "01001100101101",
                             10183 when "01001100101110",
                             10181 when "01001100101111",
                             10179 when "01001100110000",
                             10177 when "01001100110001",
                             10175 when "01001100110010",
                             10173 when "01001100110011",
                             10171 when "01001100110100",
                             10169 when "01001100110101",
                             10167 when "01001100110110",
                             10165 when "01001100110111",
                             10163 when "01001100111000",
                             10161 when "01001100111001",
                             10158 when "01001100111010",
                             10156 when "01001100111011",
                             10154 when "01001100111100",
                             10152 when "01001100111101",
                             10150 when "01001100111110",
                             10148 when "01001100111111",
                             10146 when "01001101000000",
                             10144 when "01001101000001",
                             10142 when "01001101000010",
                             10140 when "01001101000011",
                             10138 when "01001101000100",
                             10136 when "01001101000101",
                             10134 when "01001101000110",
                             10132 when "01001101000111",
                             10130 when "01001101001000",
                             10128 when "01001101001001",
                             10126 when "01001101001010",
                             10124 when "01001101001011",
                             10121 when "01001101001100",
                             10119 when "01001101001101",
                             10117 when "01001101001110",
                             10115 when "01001101001111",
                             10113 when "01001101010000",
                             10111 when "01001101010001",
                             10109 when "01001101010010",
                             10107 when "01001101010011",
                             10105 when "01001101010100",
                             10103 when "01001101010101",
                             10101 when "01001101010110",
                             10099 when "01001101010111",
                             10097 when "01001101011000",
                             10095 when "01001101011001",
                             10093 when "01001101011010",
                             10091 when "01001101011011",
                             10089 when "01001101011100",
                             10087 when "01001101011101",
                             10085 when "01001101011110",
                             10083 when "01001101011111",
                             10081 when "01001101100000",
                             10079 when "01001101100001",
                             10077 when "01001101100010",
                             10075 when "01001101100011",
                             10073 when "01001101100100",
                             10070 when "01001101100101",
                             10068 when "01001101100110",
                             10066 when "01001101100111",
                             10064 when "01001101101000",
                             10062 when "01001101101001",
                             10060 when "01001101101010",
                             10058 when "01001101101011",
                             10056 when "01001101101100",
                             10054 when "01001101101101",
                             10052 when "01001101101110",
                             10050 when "01001101101111",
                             10048 when "01001101110000",
                             10046 when "01001101110001",
                             10044 when "01001101110010",
                             10042 when "01001101110011",
                             10040 when "01001101110100",
                             10038 when "01001101110101",
                             10036 when "01001101110110",
                             10034 when "01001101110111",
                             10032 when "01001101111000",
                             10030 when "01001101111001",
                             10028 when "01001101111010",
                             10026 when "01001101111011",
                             10024 when "01001101111100",
                             10022 when "01001101111101",
                             10020 when "01001101111110",
                             10018 when "01001101111111",
                             10016 when "01001110000000",
                             10014 when "01001110000001",
                             10012 when "01001110000010",
                             10010 when "01001110000011",
                             10008 when "01001110000100",
                             10006 when "01001110000101",
                             10004 when "01001110000110",
                             10002 when "01001110000111",
                             10000 when "01001110001000",
                             9998 when "01001110001001",
                             9996 when "01001110001010",
                             9994 when "01001110001011",
                             9992 when "01001110001100",
                             9990 when "01001110001101",
                             9988 when "01001110001110",
                             9986 when "01001110001111",
                             9984 when "01001110010000",
                             9982 when "01001110010001",
                             9980 when "01001110010010",
                             9978 when "01001110010011",
                             9976 when "01001110010100",
                             9974 when "01001110010101",
                             9972 when "01001110010110",
                             9970 when "01001110010111",
                             9968 when "01001110011000",
                             9966 when "01001110011001",
                             9964 when "01001110011010",
                             9962 when "01001110011011",
                             9960 when "01001110011100",
                             9958 when "01001110011101",
                             9956 when "01001110011110",
                             9954 when "01001110011111",
                             9952 when "01001110100000",
                             9950 when "01001110100001",
                             9948 when "01001110100010",
                             9946 when "01001110100011",
                             9944 when "01001110100100",
                             9942 when "01001110100101",
                             9940 when "01001110100110",
                             9938 when "01001110100111",
                             9936 when "01001110101000",
                             9934 when "01001110101001",
                             9932 when "01001110101010",
                             9930 when "01001110101011",
                             9929 when "01001110101100",
                             9927 when "01001110101101",
                             9925 when "01001110101110",
                             9923 when "01001110101111",
                             9921 when "01001110110000",
                             9919 when "01001110110001",
                             9917 when "01001110110010",
                             9915 when "01001110110011",
                             9913 when "01001110110100",
                             9911 when "01001110110101",
                             9909 when "01001110110110",
                             9907 when "01001110110111",
                             9905 when "01001110111000",
                             9903 when "01001110111001",
                             9901 when "01001110111010",
                             9899 when "01001110111011",
                             9897 when "01001110111100",
                             9895 when "01001110111101",
                             9893 when "01001110111110",
                             9891 when "01001110111111",
                             9889 when "01001111000000",
                             9887 when "01001111000001",
                             9885 when "01001111000010",
                             9883 when "01001111000011",
                             9881 when "01001111000100",
                             9879 when "01001111000101",
                             9878 when "01001111000110",
                             9876 when "01001111000111",
                             9874 when "01001111001000",
                             9872 when "01001111001001",
                             9870 when "01001111001010",
                             9868 when "01001111001011",
                             9866 when "01001111001100",
                             9864 when "01001111001101",
                             9862 when "01001111001110",
                             9860 when "01001111001111",
                             9858 when "01001111010000",
                             9856 when "01001111010001",
                             9854 when "01001111010010",
                             9852 when "01001111010011",
                             9850 when "01001111010100",
                             9848 when "01001111010101",
                             9846 when "01001111010110",
                             9844 when "01001111010111",
                             9843 when "01001111011000",
                             9841 when "01001111011001",
                             9839 when "01001111011010",
                             9837 when "01001111011011",
                             9835 when "01001111011100",
                             9833 when "01001111011101",
                             9831 when "01001111011110",
                             9829 when "01001111011111",
                             9827 when "01001111100000",
                             9825 when "01001111100001",
                             9823 when "01001111100010",
                             9821 when "01001111100011",
                             9819 when "01001111100100",
                             9817 when "01001111100101",
                             9815 when "01001111100110",
                             9814 when "01001111100111",
                             9812 when "01001111101000",
                             9810 when "01001111101001",
                             9808 when "01001111101010",
                             9806 when "01001111101011",
                             9804 when "01001111101100",
                             9802 when "01001111101101",
                             9800 when "01001111101110",
                             9798 when "01001111101111",
                             9796 when "01001111110000",
                             9794 when "01001111110001",
                             9792 when "01001111110010",
                             9790 when "01001111110011",
                             9789 when "01001111110100",
                             9787 when "01001111110101",
                             9785 when "01001111110110",
                             9783 when "01001111110111",
                             9781 when "01001111111000",
                             9779 when "01001111111001",
                             9777 when "01001111111010",
                             9775 when "01001111111011",
                             9773 when "01001111111100",
                             9771 when "01001111111101",
                             9769 when "01001111111110",
                             9768 when "01001111111111",
                             9766 when "01010000000000",
                             9764 when "01010000000001",
                             9762 when "01010000000010",
                             9760 when "01010000000011",
                             9758 when "01010000000100",
                             9756 when "01010000000101",
                             9754 when "01010000000110",
                             9752 when "01010000000111",
                             9750 when "01010000001000",
                             9748 when "01010000001001",
                             9747 when "01010000001010",
                             9745 when "01010000001011",
                             9743 when "01010000001100",
                             9741 when "01010000001101",
                             9739 when "01010000001110",
                             9737 when "01010000001111",
                             9735 when "01010000010000",
                             9733 when "01010000010001",
                             9731 when "01010000010010",
                             9730 when "01010000010011",
                             9728 when "01010000010100",
                             9726 when "01010000010101",
                             9724 when "01010000010110",
                             9722 when "01010000010111",
                             9720 when "01010000011000",
                             9718 when "01010000011001",
                             9716 when "01010000011010",
                             9714 when "01010000011011",
                             9713 when "01010000011100",
                             9711 when "01010000011101",
                             9709 when "01010000011110",
                             9707 when "01010000011111",
                             9705 when "01010000100000",
                             9703 when "01010000100001",
                             9701 when "01010000100010",
                             9699 when "01010000100011",
                             9697 when "01010000100100",
                             9696 when "01010000100101",
                             9694 when "01010000100110",
                             9692 when "01010000100111",
                             9690 when "01010000101000",
                             9688 when "01010000101001",
                             9686 when "01010000101010",
                             9684 when "01010000101011",
                             9682 when "01010000101100",
                             9681 when "01010000101101",
                             9679 when "01010000101110",
                             9677 when "01010000101111",
                             9675 when "01010000110000",
                             9673 when "01010000110001",
                             9671 when "01010000110010",
                             9669 when "01010000110011",
                             9667 when "01010000110100",
                             9666 when "01010000110101",
                             9664 when "01010000110110",
                             9662 when "01010000110111",
                             9660 when "01010000111000",
                             9658 when "01010000111001",
                             9656 when "01010000111010",
                             9654 when "01010000111011",
                             9653 when "01010000111100",
                             9651 when "01010000111101",
                             9649 when "01010000111110",
                             9647 when "01010000111111",
                             9645 when "01010001000000",
                             9643 when "01010001000001",
                             9641 when "01010001000010",
                             9639 when "01010001000011",
                             9638 when "01010001000100",
                             9636 when "01010001000101",
                             9634 when "01010001000110",
                             9632 when "01010001000111",
                             9630 when "01010001001000",
                             9628 when "01010001001001",
                             9626 when "01010001001010",
                             9625 when "01010001001011",
                             9623 when "01010001001100",
                             9621 when "01010001001101",
                             9619 when "01010001001110",
                             9617 when "01010001001111",
                             9615 when "01010001010000",
                             9614 when "01010001010001",
                             9612 when "01010001010010",
                             9610 when "01010001010011",
                             9608 when "01010001010100",
                             9606 when "01010001010101",
                             9604 when "01010001010110",
                             9602 when "01010001010111",
                             9601 when "01010001011000",
                             9599 when "01010001011001",
                             9597 when "01010001011010",
                             9595 when "01010001011011",
                             9593 when "01010001011100",
                             9591 when "01010001011101",
                             9590 when "01010001011110",
                             9588 when "01010001011111",
                             9586 when "01010001100000",
                             9584 when "01010001100001",
                             9582 when "01010001100010",
                             9580 when "01010001100011",
                             9579 when "01010001100100",
                             9577 when "01010001100101",
                             9575 when "01010001100110",
                             9573 when "01010001100111",
                             9571 when "01010001101000",
                             9569 when "01010001101001",
                             9568 when "01010001101010",
                             9566 when "01010001101011",
                             9564 when "01010001101100",
                             9562 when "01010001101101",
                             9560 when "01010001101110",
                             9558 when "01010001101111",
                             9557 when "01010001110000",
                             9555 when "01010001110001",
                             9553 when "01010001110010",
                             9551 when "01010001110011",
                             9549 when "01010001110100",
                             9547 when "01010001110101",
                             9546 when "01010001110110",
                             9544 when "01010001110111",
                             9542 when "01010001111000",
                             9540 when "01010001111001",
                             9538 when "01010001111010",
                             9537 when "01010001111011",
                             9535 when "01010001111100",
                             9533 when "01010001111101",
                             9531 when "01010001111110",
                             9529 when "01010001111111",
                             9527 when "01010010000000",
                             9526 when "01010010000001",
                             9524 when "01010010000010",
                             9522 when "01010010000011",
                             9520 when "01010010000100",
                             9518 when "01010010000101",
                             9517 when "01010010000110",
                             9515 when "01010010000111",
                             9513 when "01010010001000",
                             9511 when "01010010001001",
                             9509 when "01010010001010",
                             9508 when "01010010001011",
                             9506 when "01010010001100",
                             9504 when "01010010001101",
                             9502 when "01010010001110",
                             9500 when "01010010001111",
                             9498 when "01010010010000",
                             9497 when "01010010010001",
                             9495 when "01010010010010",
                             9493 when "01010010010011",
                             9491 when "01010010010100",
                             9489 when "01010010010101",
                             9488 when "01010010010110",
                             9486 when "01010010010111",
                             9484 when "01010010011000",
                             9482 when "01010010011001",
                             9480 when "01010010011010",
                             9479 when "01010010011011",
                             9477 when "01010010011100",
                             9475 when "01010010011101",
                             9473 when "01010010011110",
                             9471 when "01010010011111",
                             9470 when "01010010100000",
                             9468 when "01010010100001",
                             9466 when "01010010100010",
                             9464 when "01010010100011",
                             9463 when "01010010100100",
                             9461 when "01010010100101",
                             9459 when "01010010100110",
                             9457 when "01010010100111",
                             9455 when "01010010101000",
                             9454 when "01010010101001",
                             9452 when "01010010101010",
                             9450 when "01010010101011",
                             9448 when "01010010101100",
                             9446 when "01010010101101",
                             9445 when "01010010101110",
                             9443 when "01010010101111",
                             9441 when "01010010110000",
                             9439 when "01010010110001",
                             9438 when "01010010110010",
                             9436 when "01010010110011",
                             9434 when "01010010110100",
                             9432 when "01010010110101",
                             9430 when "01010010110110",
                             9429 when "01010010110111",
                             9427 when "01010010111000",
                             9425 when "01010010111001",
                             9423 when "01010010111010",
                             9422 when "01010010111011",
                             9420 when "01010010111100",
                             9418 when "01010010111101",
                             9416 when "01010010111110",
                             9414 when "01010010111111",
                             9413 when "01010011000000",
                             9411 when "01010011000001",
                             9409 when "01010011000010",
                             9407 when "01010011000011",
                             9406 when "01010011000100",
                             9404 when "01010011000101",
                             9402 when "01010011000110",
                             9400 when "01010011000111",
                             9398 when "01010011001000",
                             9397 when "01010011001001",
                             9395 when "01010011001010",
                             9393 when "01010011001011",
                             9391 when "01010011001100",
                             9390 when "01010011001101",
                             9388 when "01010011001110",
                             9386 when "01010011001111",
                             9384 when "01010011010000",
                             9383 when "01010011010001",
                             9381 when "01010011010010",
                             9379 when "01010011010011",
                             9377 when "01010011010100",
                             9376 when "01010011010101",
                             9374 when "01010011010110",
                             9372 when "01010011010111",
                             9370 when "01010011011000",
                             9369 when "01010011011001",
                             9367 when "01010011011010",
                             9365 when "01010011011011",
                             9363 when "01010011011100",
                             9362 when "01010011011101",
                             9360 when "01010011011110",
                             9358 when "01010011011111",
                             9356 when "01010011100000",
                             9355 when "01010011100001",
                             9353 when "01010011100010",
                             9351 when "01010011100011",
                             9349 when "01010011100100",
                             9348 when "01010011100101",
                             9346 when "01010011100110",
                             9344 when "01010011100111",
                             9342 when "01010011101000",
                             9341 when "01010011101001",
                             9339 when "01010011101010",
                             9337 when "01010011101011",
                             9335 when "01010011101100",
                             9334 when "01010011101101",
                             9332 when "01010011101110",
                             9330 when "01010011101111",
                             9328 when "01010011110000",
                             9327 when "01010011110001",
                             9325 when "01010011110010",
                             9323 when "01010011110011",
                             9321 when "01010011110100",
                             9320 when "01010011110101",
                             9318 when "01010011110110",
                             9316 when "01010011110111",
                             9314 when "01010011111000",
                             9313 when "01010011111001",
                             9311 when "01010011111010",
                             9309 when "01010011111011",
                             9308 when "01010011111100",
                             9306 when "01010011111101",
                             9304 when "01010011111110",
                             9302 when "01010011111111",
                             9301 when "01010100000000",
                             9299 when "01010100000001",
                             9297 when "01010100000010",
                             9295 when "01010100000011",
                             9294 when "01010100000100",
                             9292 when "01010100000101",
                             9290 when "01010100000110",
                             9289 when "01010100000111",
                             9287 when "01010100001000",
                             9285 when "01010100001001",
                             9283 when "01010100001010",
                             9282 when "01010100001011",
                             9280 when "01010100001100",
                             9278 when "01010100001101",
                             9276 when "01010100001110",
                             9275 when "01010100001111",
                             9273 when "01010100010000",
                             9271 when "01010100010001",
                             9270 when "01010100010010",
                             9268 when "01010100010011",
                             9266 when "01010100010100",
                             9264 when "01010100010101",
                             9263 when "01010100010110",
                             9261 when "01010100010111",
                             9259 when "01010100011000",
                             9258 when "01010100011001",
                             9256 when "01010100011010",
                             9254 when "01010100011011",
                             9252 when "01010100011100",
                             9251 when "01010100011101",
                             9249 when "01010100011110",
                             9247 when "01010100011111",
                             9246 when "01010100100000",
                             9244 when "01010100100001",
                             9242 when "01010100100010",
                             9240 when "01010100100011",
                             9239 when "01010100100100",
                             9237 when "01010100100101",
                             9235 when "01010100100110",
                             9234 when "01010100100111",
                             9232 when "01010100101000",
                             9230 when "01010100101001",
                             9228 when "01010100101010",
                             9227 when "01010100101011",
                             9225 when "01010100101100",
                             9223 when "01010100101101",
                             9222 when "01010100101110",
                             9220 when "01010100101111",
                             9218 when "01010100110000",
                             9217 when "01010100110001",
                             9215 when "01010100110010",
                             9213 when "01010100110011",
                             9211 when "01010100110100",
                             9210 when "01010100110101",
                             9208 when "01010100110110",
                             9206 when "01010100110111",
                             9205 when "01010100111000",
                             9203 when "01010100111001",
                             9201 when "01010100111010",
                             9200 when "01010100111011",
                             9198 when "01010100111100",
                             9196 when "01010100111101",
                             9195 when "01010100111110",
                             9193 when "01010100111111",
                             9191 when "01010101000000",
                             9189 when "01010101000001",
                             9188 when "01010101000010",
                             9186 when "01010101000011",
                             9184 when "01010101000100",
                             9183 when "01010101000101",
                             9181 when "01010101000110",
                             9179 when "01010101000111",
                             9178 when "01010101001000",
                             9176 when "01010101001001",
                             9174 when "01010101001010",
                             9173 when "01010101001011",
                             9171 when "01010101001100",
                             9169 when "01010101001101",
                             9168 when "01010101001110",
                             9166 when "01010101001111",
                             9164 when "01010101010000",
                             9163 when "01010101010001",
                             9161 when "01010101010010",
                             9159 when "01010101010011",
                             9158 when "01010101010100",
                             9156 when "01010101010101",
                             9154 when "01010101010110",
                             9152 when "01010101010111",
                             9151 when "01010101011000",
                             9149 when "01010101011001",
                             9147 when "01010101011010",
                             9146 when "01010101011011",
                             9144 when "01010101011100",
                             9142 when "01010101011101",
                             9141 when "01010101011110",
                             9139 when "01010101011111",
                             9137 when "01010101100000",
                             9136 when "01010101100001",
                             9134 when "01010101100010",
                             9132 when "01010101100011",
                             9131 when "01010101100100",
                             9129 when "01010101100101",
                             9127 when "01010101100110",
                             9126 when "01010101100111",
                             9124 when "01010101101000",
                             9122 when "01010101101001",
                             9121 when "01010101101010",
                             9119 when "01010101101011",
                             9117 when "01010101101100",
                             9116 when "01010101101101",
                             9114 when "01010101101110",
                             9112 when "01010101101111",
                             9111 when "01010101110000",
                             9109 when "01010101110001",
                             9107 when "01010101110010",
                             9106 when "01010101110011",
                             9104 when "01010101110100",
                             9102 when "01010101110101",
                             9101 when "01010101110110",
                             9099 when "01010101110111",
                             9098 when "01010101111000",
                             9096 when "01010101111001",
                             9094 when "01010101111010",
                             9093 when "01010101111011",
                             9091 when "01010101111100",
                             9089 when "01010101111101",
                             9088 when "01010101111110",
                             9086 when "01010101111111",
                             9084 when "01010110000000",
                             9083 when "01010110000001",
                             9081 when "01010110000010",
                             9079 when "01010110000011",
                             9078 when "01010110000100",
                             9076 when "01010110000101",
                             9074 when "01010110000110",
                             9073 when "01010110000111",
                             9071 when "01010110001000",
                             9069 when "01010110001001",
                             9068 when "01010110001010",
                             9066 when "01010110001011",
                             9065 when "01010110001100",
                             9063 when "01010110001101",
                             9061 when "01010110001110",
                             9060 when "01010110001111",
                             9058 when "01010110010000",
                             9056 when "01010110010001",
                             9055 when "01010110010010",
                             9053 when "01010110010011",
                             9051 when "01010110010100",
                             9050 when "01010110010101",
                             9048 when "01010110010110",
                             9046 when "01010110010111",
                             9045 when "01010110011000",
                             9043 when "01010110011001",
                             9042 when "01010110011010",
                             9040 when "01010110011011",
                             9038 when "01010110011100",
                             9037 when "01010110011101",
                             9035 when "01010110011110",
                             9033 when "01010110011111",
                             9032 when "01010110100000",
                             9030 when "01010110100001",
                             9029 when "01010110100010",
                             9027 when "01010110100011",
                             9025 when "01010110100100",
                             9024 when "01010110100101",
                             9022 when "01010110100110",
                             9020 when "01010110100111",
                             9019 when "01010110101000",
                             9017 when "01010110101001",
                             9016 when "01010110101010",
                             9014 when "01010110101011",
                             9012 when "01010110101100",
                             9011 when "01010110101101",
                             9009 when "01010110101110",
                             9007 when "01010110101111",
                             9006 when "01010110110000",
                             9004 when "01010110110001",
                             9003 when "01010110110010",
                             9001 when "01010110110011",
                             8999 when "01010110110100",
                             8998 when "01010110110101",
                             8996 when "01010110110110",
                             8994 when "01010110110111",
                             8993 when "01010110111000",
                             8991 when "01010110111001",
                             8990 when "01010110111010",
                             8988 when "01010110111011",
                             8986 when "01010110111100",
                             8985 when "01010110111101",
                             8983 when "01010110111110",
                             8981 when "01010110111111",
                             8980 when "01010111000000",
                             8978 when "01010111000001",
                             8977 when "01010111000010",
                             8975 when "01010111000011",
                             8973 when "01010111000100",
                             8972 when "01010111000101",
                             8970 when "01010111000110",
                             8969 when "01010111000111",
                             8967 when "01010111001000",
                             8965 when "01010111001001",
                             8964 when "01010111001010",
                             8962 when "01010111001011",
                             8961 when "01010111001100",
                             8959 when "01010111001101",
                             8957 when "01010111001110",
                             8956 when "01010111001111",
                             8954 when "01010111010000",
                             8953 when "01010111010001",
                             8951 when "01010111010010",
                             8949 when "01010111010011",
                             8948 when "01010111010100",
                             8946 when "01010111010101",
                             8945 when "01010111010110",
                             8943 when "01010111010111",
                             8941 when "01010111011000",
                             8940 when "01010111011001",
                             8938 when "01010111011010",
                             8937 when "01010111011011",
                             8935 when "01010111011100",
                             8933 when "01010111011101",
                             8932 when "01010111011110",
                             8930 when "01010111011111",
                             8929 when "01010111100000",
                             8927 when "01010111100001",
                             8925 when "01010111100010",
                             8924 when "01010111100011",
                             8922 when "01010111100100",
                             8921 when "01010111100101",
                             8919 when "01010111100110",
                             8917 when "01010111100111",
                             8916 when "01010111101000",
                             8914 when "01010111101001",
                             8913 when "01010111101010",
                             8911 when "01010111101011",
                             8909 when "01010111101100",
                             8908 when "01010111101101",
                             8906 when "01010111101110",
                             8905 when "01010111101111",
                             8903 when "01010111110000",
                             8902 when "01010111110001",
                             8900 when "01010111110010",
                             8898 when "01010111110011",
                             8897 when "01010111110100",
                             8895 when "01010111110101",
                             8894 when "01010111110110",
                             8892 when "01010111110111",
                             8890 when "01010111111000",
                             8889 when "01010111111001",
                             8887 when "01010111111010",
                             8886 when "01010111111011",
                             8884 when "01010111111100",
                             8883 when "01010111111101",
                             8881 when "01010111111110",
                             8879 when "01010111111111",
                             8878 when "01011000000000",
                             8876 when "01011000000001",
                             8875 when "01011000000010",
                             8873 when "01011000000011",
                             8872 when "01011000000100",
                             8870 when "01011000000101",
                             8868 when "01011000000110",
                             8867 when "01011000000111",
                             8865 when "01011000001000",
                             8864 when "01011000001001",
                             8862 when "01011000001010",
                             8861 when "01011000001011",
                             8859 when "01011000001100",
                             8857 when "01011000001101",
                             8856 when "01011000001110",
                             8854 when "01011000001111",
                             8853 when "01011000010000",
                             8851 when "01011000010001",
                             8850 when "01011000010010",
                             8848 when "01011000010011",
                             8846 when "01011000010100",
                             8845 when "01011000010101",
                             8843 when "01011000010110",
                             8842 when "01011000010111",
                             8840 when "01011000011000",
                             8839 when "01011000011001",
                             8837 when "01011000011010",
                             8835 when "01011000011011",
                             8834 when "01011000011100",
                             8832 when "01011000011101",
                             8831 when "01011000011110",
                             8829 when "01011000011111",
                             8828 when "01011000100000",
                             8826 when "01011000100001",
                             8825 when "01011000100010",
                             8823 when "01011000100011",
                             8821 when "01011000100100",
                             8820 when "01011000100101",
                             8818 when "01011000100110",
                             8817 when "01011000100111",
                             8815 when "01011000101000",
                             8814 when "01011000101001",
                             8812 when "01011000101010",
                             8811 when "01011000101011",
                             8809 when "01011000101100",
                             8807 when "01011000101101",
                             8806 when "01011000101110",
                             8804 when "01011000101111",
                             8803 when "01011000110000",
                             8801 when "01011000110001",
                             8800 when "01011000110010",
                             8798 when "01011000110011",
                             8797 when "01011000110100",
                             8795 when "01011000110101",
                             8794 when "01011000110110",
                             8792 when "01011000110111",
                             8790 when "01011000111000",
                             8789 when "01011000111001",
                             8787 when "01011000111010",
                             8786 when "01011000111011",
                             8784 when "01011000111100",
                             8783 when "01011000111101",
                             8781 when "01011000111110",
                             8780 when "01011000111111",
                             8778 when "01011001000000",
                             8777 when "01011001000001",
                             8775 when "01011001000010",
                             8773 when "01011001000011",
                             8772 when "01011001000100",
                             8770 when "01011001000101",
                             8769 when "01011001000110",
                             8767 when "01011001000111",
                             8766 when "01011001001000",
                             8764 when "01011001001001",
                             8763 when "01011001001010",
                             8761 when "01011001001011",
                             8760 when "01011001001100",
                             8758 when "01011001001101",
                             8757 when "01011001001110",
                             8755 when "01011001001111",
                             8754 when "01011001010000",
                             8752 when "01011001010001",
                             8750 when "01011001010010",
                             8749 when "01011001010011",
                             8747 when "01011001010100",
                             8746 when "01011001010101",
                             8744 when "01011001010110",
                             8743 when "01011001010111",
                             8741 when "01011001011000",
                             8740 when "01011001011001",
                             8738 when "01011001011010",
                             8737 when "01011001011011",
                             8735 when "01011001011100",
                             8734 when "01011001011101",
                             8732 when "01011001011110",
                             8731 when "01011001011111",
                             8729 when "01011001100000",
                             8728 when "01011001100001",
                             8726 when "01011001100010",
                             8724 when "01011001100011",
                             8723 when "01011001100100",
                             8721 when "01011001100101",
                             8720 when "01011001100110",
                             8718 when "01011001100111",
                             8717 when "01011001101000",
                             8715 when "01011001101001",
                             8714 when "01011001101010",
                             8712 when "01011001101011",
                             8711 when "01011001101100",
                             8709 when "01011001101101",
                             8708 when "01011001101110",
                             8706 when "01011001101111",
                             8705 when "01011001110000",
                             8703 when "01011001110001",
                             8702 when "01011001110010",
                             8700 when "01011001110011",
                             8699 when "01011001110100",
                             8697 when "01011001110101",
                             8696 when "01011001110110",
                             8694 when "01011001110111",
                             8693 when "01011001111000",
                             8691 when "01011001111001",
                             8690 when "01011001111010",
                             8688 when "01011001111011",
                             8687 when "01011001111100",
                             8685 when "01011001111101",
                             8684 when "01011001111110",
                             8682 when "01011001111111",
                             8681 when "01011010000000",
                             8679 when "01011010000001",
                             8678 when "01011010000010",
                             8676 when "01011010000011",
                             8675 when "01011010000100",
                             8673 when "01011010000101",
                             8672 when "01011010000110",
                             8670 when "01011010000111",
                             8669 when "01011010001000",
                             8667 when "01011010001001",
                             8666 when "01011010001010",
                             8664 when "01011010001011",
                             8663 when "01011010001100",
                             8661 when "01011010001101",
                             8660 when "01011010001110",
                             8658 when "01011010001111",
                             8657 when "01011010010000",
                             8655 when "01011010010001",
                             8654 when "01011010010010",
                             8652 when "01011010010011",
                             8651 when "01011010010100",
                             8649 when "01011010010101",
                             8648 when "01011010010110",
                             8646 when "01011010010111",
                             8645 when "01011010011000",
                             8643 when "01011010011001",
                             8642 when "01011010011010",
                             8640 when "01011010011011",
                             8639 when "01011010011100",
                             8637 when "01011010011101",
                             8636 when "01011010011110",
                             8634 when "01011010011111",
                             8633 when "01011010100000",
                             8631 when "01011010100001",
                             8630 when "01011010100010",
                             8628 when "01011010100011",
                             8627 when "01011010100100",
                             8625 when "01011010100101",
                             8624 when "01011010100110",
                             8622 when "01011010100111",
                             8621 when "01011010101000",
                             8619 when "01011010101001",
                             8618 when "01011010101010",
                             8616 when "01011010101011",
                             8615 when "01011010101100",
                             8613 when "01011010101101",
                             8612 when "01011010101110",
                             8610 when "01011010101111",
                             8609 when "01011010110000",
                             8607 when "01011010110001",
                             8606 when "01011010110010",
                             8604 when "01011010110011",
                             8603 when "01011010110100",
                             8601 when "01011010110101",
                             8600 when "01011010110110",
                             8598 when "01011010110111",
                             8597 when "01011010111000",
                             8595 when "01011010111001",
                             8594 when "01011010111010",
                             8593 when "01011010111011",
                             8591 when "01011010111100",
                             8590 when "01011010111101",
                             8588 when "01011010111110",
                             8587 when "01011010111111",
                             8585 when "01011011000000",
                             8584 when "01011011000001",
                             8582 when "01011011000010",
                             8581 when "01011011000011",
                             8579 when "01011011000100",
                             8578 when "01011011000101",
                             8576 when "01011011000110",
                             8575 when "01011011000111",
                             8573 when "01011011001000",
                             8572 when "01011011001001",
                             8570 when "01011011001010",
                             8569 when "01011011001011",
                             8568 when "01011011001100",
                             8566 when "01011011001101",
                             8565 when "01011011001110",
                             8563 when "01011011001111",
                             8562 when "01011011010000",
                             8560 when "01011011010001",
                             8559 when "01011011010010",
                             8557 when "01011011010011",
                             8556 when "01011011010100",
                             8554 when "01011011010101",
                             8553 when "01011011010110",
                             8551 when "01011011010111",
                             8550 when "01011011011000",
                             8548 when "01011011011001",
                             8547 when "01011011011010",
                             8546 when "01011011011011",
                             8544 when "01011011011100",
                             8543 when "01011011011101",
                             8541 when "01011011011110",
                             8540 when "01011011011111",
                             8538 when "01011011100000",
                             8537 when "01011011100001",
                             8535 when "01011011100010",
                             8534 when "01011011100011",
                             8532 when "01011011100100",
                             8531 when "01011011100101",
                             8530 when "01011011100110",
                             8528 when "01011011100111",
                             8527 when "01011011101000",
                             8525 when "01011011101001",
                             8524 when "01011011101010",
                             8522 when "01011011101011",
                             8521 when "01011011101100",
                             8519 when "01011011101101",
                             8518 when "01011011101110",
                             8516 when "01011011101111",
                             8515 when "01011011110000",
                             8514 when "01011011110001",
                             8512 when "01011011110010",
                             8511 when "01011011110011",
                             8509 when "01011011110100",
                             8508 when "01011011110101",
                             8506 when "01011011110110",
                             8505 when "01011011110111",
                             8503 when "01011011111000",
                             8502 when "01011011111001",
                             8501 when "01011011111010",
                             8499 when "01011011111011",
                             8498 when "01011011111100",
                             8496 when "01011011111101",
                             8495 when "01011011111110",
                             8493 when "01011011111111",
                             8492 when "01011100000000",
                             8490 when "01011100000001",
                             8489 when "01011100000010",
                             8488 when "01011100000011",
                             8486 when "01011100000100",
                             8485 when "01011100000101",
                             8483 when "01011100000110",
                             8482 when "01011100000111",
                             8480 when "01011100001000",
                             8479 when "01011100001001",
                             8477 when "01011100001010",
                             8476 when "01011100001011",
                             8475 when "01011100001100",
                             8473 when "01011100001101",
                             8472 when "01011100001110",
                             8470 when "01011100001111",
                             8469 when "01011100010000",
                             8467 when "01011100010001",
                             8466 when "01011100010010",
                             8465 when "01011100010011",
                             8463 when "01011100010100",
                             8462 when "01011100010101",
                             8460 when "01011100010110",
                             8459 when "01011100010111",
                             8457 when "01011100011000",
                             8456 when "01011100011001",
                             8455 when "01011100011010",
                             8453 when "01011100011011",
                             8452 when "01011100011100",
                             8450 when "01011100011101",
                             8449 when "01011100011110",
                             8447 when "01011100011111",
                             8446 when "01011100100000",
                             8445 when "01011100100001",
                             8443 when "01011100100010",
                             8442 when "01011100100011",
                             8440 when "01011100100100",
                             8439 when "01011100100101",
                             8437 when "01011100100110",
                             8436 when "01011100100111",
                             8435 when "01011100101000",
                             8433 when "01011100101001",
                             8432 when "01011100101010",
                             8430 when "01011100101011",
                             8429 when "01011100101100",
                             8427 when "01011100101101",
                             8426 when "01011100101110",
                             8425 when "01011100101111",
                             8423 when "01011100110000",
                             8422 when "01011100110001",
                             8420 when "01011100110010",
                             8419 when "01011100110011",
                             8418 when "01011100110100",
                             8416 when "01011100110101",
                             8415 when "01011100110110",
                             8413 when "01011100110111",
                             8412 when "01011100111000",
                             8410 when "01011100111001",
                             8409 when "01011100111010",
                             8408 when "01011100111011",
                             8406 when "01011100111100",
                             8405 when "01011100111101",
                             8403 when "01011100111110",
                             8402 when "01011100111111",
                             8401 when "01011101000000",
                             8399 when "01011101000001",
                             8398 when "01011101000010",
                             8396 when "01011101000011",
                             8395 when "01011101000100",
                             8393 when "01011101000101",
                             8392 when "01011101000110",
                             8391 when "01011101000111",
                             8389 when "01011101001000",
                             8388 when "01011101001001",
                             8386 when "01011101001010",
                             8385 when "01011101001011",
                             8384 when "01011101001100",
                             8382 when "01011101001101",
                             8381 when "01011101001110",
                             8379 when "01011101001111",
                             8378 when "01011101010000",
                             8377 when "01011101010001",
                             8375 when "01011101010010",
                             8374 when "01011101010011",
                             8372 when "01011101010100",
                             8371 when "01011101010101",
                             8370 when "01011101010110",
                             8368 when "01011101010111",
                             8367 when "01011101011000",
                             8365 when "01011101011001",
                             8364 when "01011101011010",
                             8363 when "01011101011011",
                             8361 when "01011101011100",
                             8360 when "01011101011101",
                             8358 when "01011101011110",
                             8357 when "01011101011111",
                             8356 when "01011101100000",
                             8354 when "01011101100001",
                             8353 when "01011101100010",
                             8351 when "01011101100011",
                             8350 when "01011101100100",
                             8349 when "01011101100101",
                             8347 when "01011101100110",
                             8346 when "01011101100111",
                             8344 when "01011101101000",
                             8343 when "01011101101001",
                             8342 when "01011101101010",
                             8340 when "01011101101011",
                             8339 when "01011101101100",
                             8338 when "01011101101101",
                             8336 when "01011101101110",
                             8335 when "01011101101111",
                             8333 when "01011101110000",
                             8332 when "01011101110001",
                             8331 when "01011101110010",
                             8329 when "01011101110011",
                             8328 when "01011101110100",
                             8326 when "01011101110101",
                             8325 when "01011101110110",
                             8324 when "01011101110111",
                             8322 when "01011101111000",
                             8321 when "01011101111001",
                             8319 when "01011101111010",
                             8318 when "01011101111011",
                             8317 when "01011101111100",
                             8315 when "01011101111101",
                             8314 when "01011101111110",
                             8313 when "01011101111111",
                             8311 when "01011110000000",
                             8310 when "01011110000001",
                             8308 when "01011110000010",
                             8307 when "01011110000011",
                             8306 when "01011110000100",
                             8304 when "01011110000101",
                             8303 when "01011110000110",
                             8302 when "01011110000111",
                             8300 when "01011110001000",
                             8299 when "01011110001001",
                             8297 when "01011110001010",
                             8296 when "01011110001011",
                             8295 when "01011110001100",
                             8293 when "01011110001101",
                             8292 when "01011110001110",
                             8290 when "01011110001111",
                             8289 when "01011110010000",
                             8288 when "01011110010001",
                             8286 when "01011110010010",
                             8285 when "01011110010011",
                             8284 when "01011110010100",
                             8282 when "01011110010101",
                             8281 when "01011110010110",
                             8280 when "01011110010111",
                             8278 when "01011110011000",
                             8277 when "01011110011001",
                             8275 when "01011110011010",
                             8274 when "01011110011011",
                             8273 when "01011110011100",
                             8271 when "01011110011101",
                             8270 when "01011110011110",
                             8269 when "01011110011111",
                             8267 when "01011110100000",
                             8266 when "01011110100001",
                             8264 when "01011110100010",
                             8263 when "01011110100011",
                             8262 when "01011110100100",
                             8260 when "01011110100101",
                             8259 when "01011110100110",
                             8258 when "01011110100111",
                             8256 when "01011110101000",
                             8255 when "01011110101001",
                             8254 when "01011110101010",
                             8252 when "01011110101011",
                             8251 when "01011110101100",
                             8249 when "01011110101101",
                             8248 when "01011110101110",
                             8247 when "01011110101111",
                             8245 when "01011110110000",
                             8244 when "01011110110001",
                             8243 when "01011110110010",
                             8241 when "01011110110011",
                             8240 when "01011110110100",
                             8239 when "01011110110101",
                             8237 when "01011110110110",
                             8236 when "01011110110111",
                             8235 when "01011110111000",
                             8233 when "01011110111001",
                             8232 when "01011110111010",
                             8230 when "01011110111011",
                             8229 when "01011110111100",
                             8228 when "01011110111101",
                             8226 when "01011110111110",
                             8225 when "01011110111111",
                             8224 when "01011111000000",
                             8222 when "01011111000001",
                             8221 when "01011111000010",
                             8220 when "01011111000011",
                             8218 when "01011111000100",
                             8217 when "01011111000101",
                             8216 when "01011111000110",
                             8214 when "01011111000111",
                             8213 when "01011111001000",
                             8212 when "01011111001001",
                             8210 when "01011111001010",
                             8209 when "01011111001011",
                             8207 when "01011111001100",
                             8206 when "01011111001101",
                             8205 when "01011111001110",
                             8203 when "01011111001111",
                             8202 when "01011111010000",
                             8201 when "01011111010001",
                             8199 when "01011111010010",
                             8198 when "01011111010011",
                             8197 when "01011111010100",
                             8195 when "01011111010101",
                             8194 when "01011111010110",
                             8193 when "01011111010111",
                             8191 when "01011111011000",
                             8190 when "01011111011001",
                             8189 when "01011111011010",
                             8187 when "01011111011011",
                             8186 when "01011111011100",
                             8185 when "01011111011101",
                             8183 when "01011111011110",
                             8182 when "01011111011111",
                             8181 when "01011111100000",
                             8179 when "01011111100001",
                             8178 when "01011111100010",
                             8177 when "01011111100011",
                             8175 when "01011111100100",
                             8174 when "01011111100101",
                             8173 when "01011111100110",
                             8171 when "01011111100111",
                             8170 when "01011111101000",
                             8169 when "01011111101001",
                             8167 when "01011111101010",
                             8166 when "01011111101011",
                             8165 when "01011111101100",
                             8163 when "01011111101101",
                             8162 when "01011111101110",
                             8161 when "01011111101111",
                             8159 when "01011111110000",
                             8158 when "01011111110001",
                             8157 when "01011111110010",
                             8155 when "01011111110011",
                             8154 when "01011111110100",
                             8153 when "01011111110101",
                             8151 when "01011111110110",
                             8150 when "01011111110111",
                             8149 when "01011111111000",
                             8147 when "01011111111001",
                             8146 when "01011111111010",
                             8145 when "01011111111011",
                             8143 when "01011111111100",
                             8142 when "01011111111101",
                             8141 when "01011111111110",
                             8139 when "01011111111111",
                             8138 when "01100000000000",
                             8137 when "01100000000001",
                             8135 when "01100000000010",
                             8134 when "01100000000011",
                             8133 when "01100000000100",
                             8131 when "01100000000101",
                             8130 when "01100000000110",
                             8129 when "01100000000111",
                             8127 when "01100000001000",
                             8126 when "01100000001001",
                             8125 when "01100000001010",
                             8123 when "01100000001011",
                             8122 when "01100000001100",
                             8121 when "01100000001101",
                             8120 when "01100000001110",
                             8118 when "01100000001111",
                             8117 when "01100000010000",
                             8116 when "01100000010001",
                             8114 when "01100000010010",
                             8113 when "01100000010011",
                             8112 when "01100000010100",
                             8110 when "01100000010101",
                             8109 when "01100000010110",
                             8108 when "01100000010111",
                             8106 when "01100000011000",
                             8105 when "01100000011001",
                             8104 when "01100000011010",
                             8102 when "01100000011011",
                             8101 when "01100000011100",
                             8100 when "01100000011101",
                             8098 when "01100000011110",
                             8097 when "01100000011111",
                             8096 when "01100000100000",
                             8095 when "01100000100001",
                             8093 when "01100000100010",
                             8092 when "01100000100011",
                             8091 when "01100000100100",
                             8089 when "01100000100101",
                             8088 when "01100000100110",
                             8087 when "01100000100111",
                             8085 when "01100000101000",
                             8084 when "01100000101001",
                             8083 when "01100000101010",
                             8081 when "01100000101011",
                             8080 when "01100000101100",
                             8079 when "01100000101101",
                             8078 when "01100000101110",
                             8076 when "01100000101111",
                             8075 when "01100000110000",
                             8074 when "01100000110001",
                             8072 when "01100000110010",
                             8071 when "01100000110011",
                             8070 when "01100000110100",
                             8068 when "01100000110101",
                             8067 when "01100000110110",
                             8066 when "01100000110111",
                             8065 when "01100000111000",
                             8063 when "01100000111001",
                             8062 when "01100000111010",
                             8061 when "01100000111011",
                             8059 when "01100000111100",
                             8058 when "01100000111101",
                             8057 when "01100000111110",
                             8055 when "01100000111111",
                             8054 when "01100001000000",
                             8053 when "01100001000001",
                             8052 when "01100001000010",
                             8050 when "01100001000011",
                             8049 when "01100001000100",
                             8048 when "01100001000101",
                             8046 when "01100001000110",
                             8045 when "01100001000111",
                             8044 when "01100001001000",
                             8042 when "01100001001001",
                             8041 when "01100001001010",
                             8040 when "01100001001011",
                             8039 when "01100001001100",
                             8037 when "01100001001101",
                             8036 when "01100001001110",
                             8035 when "01100001001111",
                             8033 when "01100001010000",
                             8032 when "01100001010001",
                             8031 when "01100001010010",
                             8030 when "01100001010011",
                             8028 when "01100001010100",
                             8027 when "01100001010101",
                             8026 when "01100001010110",
                             8024 when "01100001010111",
                             8023 when "01100001011000",
                             8022 when "01100001011001",
                             8021 when "01100001011010",
                             8019 when "01100001011011",
                             8018 when "01100001011100",
                             8017 when "01100001011101",
                             8015 when "01100001011110",
                             8014 when "01100001011111",
                             8013 when "01100001100000",
                             8012 when "01100001100001",
                             8010 when "01100001100010",
                             8009 when "01100001100011",
                             8008 when "01100001100100",
                             8006 when "01100001100101",
                             8005 when "01100001100110",
                             8004 when "01100001100111",
                             8003 when "01100001101000",
                             8001 when "01100001101001",
                             8000 when "01100001101010",
                             7999 when "01100001101011",
                             7997 when "01100001101100",
                             7996 when "01100001101101",
                             7995 when "01100001101110",
                             7994 when "01100001101111",
                             7992 when "01100001110000",
                             7991 when "01100001110001",
                             7990 when "01100001110010",
                             7988 when "01100001110011",
                             7987 when "01100001110100",
                             7986 when "01100001110101",
                             7985 when "01100001110110",
                             7983 when "01100001110111",
                             7982 when "01100001111000",
                             7981 when "01100001111001",
                             7980 when "01100001111010",
                             7978 when "01100001111011",
                             7977 when "01100001111100",
                             7976 when "01100001111101",
                             7974 when "01100001111110",
                             7973 when "01100001111111",
                             7972 when "01100010000000",
                             7971 when "01100010000001",
                             7969 when "01100010000010",
                             7968 when "01100010000011",
                             7967 when "01100010000100",
                             7966 when "01100010000101",
                             7964 when "01100010000110",
                             7963 when "01100010000111",
                             7962 when "01100010001000",
                             7961 when "01100010001001",
                             7959 when "01100010001010",
                             7958 when "01100010001011",
                             7957 when "01100010001100",
                             7955 when "01100010001101",
                             7954 when "01100010001110",
                             7953 when "01100010001111",
                             7952 when "01100010010000",
                             7950 when "01100010010001",
                             7949 when "01100010010010",
                             7948 when "01100010010011",
                             7947 when "01100010010100",
                             7945 when "01100010010101",
                             7944 when "01100010010110",
                             7943 when "01100010010111",
                             7942 when "01100010011000",
                             7940 when "01100010011001",
                             7939 when "01100010011010",
                             7938 when "01100010011011",
                             7937 when "01100010011100",
                             7935 when "01100010011101",
                             7934 when "01100010011110",
                             7933 when "01100010011111",
                             7931 when "01100010100000",
                             7930 when "01100010100001",
                             7929 when "01100010100010",
                             7928 when "01100010100011",
                             7926 when "01100010100100",
                             7925 when "01100010100101",
                             7924 when "01100010100110",
                             7923 when "01100010100111",
                             7921 when "01100010101000",
                             7920 when "01100010101001",
                             7919 when "01100010101010",
                             7918 when "01100010101011",
                             7916 when "01100010101100",
                             7915 when "01100010101101",
                             7914 when "01100010101110",
                             7913 when "01100010101111",
                             7911 when "01100010110000",
                             7910 when "01100010110001",
                             7909 when "01100010110010",
                             7908 when "01100010110011",
                             7906 when "01100010110100",
                             7905 when "01100010110101",
                             7904 when "01100010110110",
                             7903 when "01100010110111",
                             7901 when "01100010111000",
                             7900 when "01100010111001",
                             7899 when "01100010111010",
                             7898 when "01100010111011",
                             7896 when "01100010111100",
                             7895 when "01100010111101",
                             7894 when "01100010111110",
                             7893 when "01100010111111",
                             7891 when "01100011000000",
                             7890 when "01100011000001",
                             7889 when "01100011000010",
                             7888 when "01100011000011",
                             7886 when "01100011000100",
                             7885 when "01100011000101",
                             7884 when "01100011000110",
                             7883 when "01100011000111",
                             7881 when "01100011001000",
                             7880 when "01100011001001",
                             7879 when "01100011001010",
                             7878 when "01100011001011",
                             7876 when "01100011001100",
                             7875 when "01100011001101",
                             7874 when "01100011001110",
                             7873 when "01100011001111",
                             7872 when "01100011010000",
                             7870 when "01100011010001",
                             7869 when "01100011010010",
                             7868 when "01100011010011",
                             7867 when "01100011010100",
                             7865 when "01100011010101",
                             7864 when "01100011010110",
                             7863 when "01100011010111",
                             7862 when "01100011011000",
                             7860 when "01100011011001",
                             7859 when "01100011011010",
                             7858 when "01100011011011",
                             7857 when "01100011011100",
                             7855 when "01100011011101",
                             7854 when "01100011011110",
                             7853 when "01100011011111",
                             7852 when "01100011100000",
                             7851 when "01100011100001",
                             7849 when "01100011100010",
                             7848 when "01100011100011",
                             7847 when "01100011100100",
                             7846 when "01100011100101",
                             7844 when "01100011100110",
                             7843 when "01100011100111",
                             7842 when "01100011101000",
                             7841 when "01100011101001",
                             7839 when "01100011101010",
                             7838 when "01100011101011",
                             7837 when "01100011101100",
                             7836 when "01100011101101",
                             7835 when "01100011101110",
                             7833 when "01100011101111",
                             7832 when "01100011110000",
                             7831 when "01100011110001",
                             7830 when "01100011110010",
                             7828 when "01100011110011",
                             7827 when "01100011110100",
                             7826 when "01100011110101",
                             7825 when "01100011110110",
                             7824 when "01100011110111",
                             7822 when "01100011111000",
                             7821 when "01100011111001",
                             7820 when "01100011111010",
                             7819 when "01100011111011",
                             7817 when "01100011111100",
                             7816 when "01100011111101",
                             7815 when "01100011111110",
                             7814 when "01100011111111",
                             7813 when "01100100000000",
                             7811 when "01100100000001",
                             7810 when "01100100000010",
                             7809 when "01100100000011",
                             7808 when "01100100000100",
                             7806 when "01100100000101",
                             7805 when "01100100000110",
                             7804 when "01100100000111",
                             7803 when "01100100001000",
                             7802 when "01100100001001",
                             7800 when "01100100001010",
                             7799 when "01100100001011",
                             7798 when "01100100001100",
                             7797 when "01100100001101",
                             7795 when "01100100001110",
                             7794 when "01100100001111",
                             7793 when "01100100010000",
                             7792 when "01100100010001",
                             7791 when "01100100010010",
                             7789 when "01100100010011",
                             7788 when "01100100010100",
                             7787 when "01100100010101",
                             7786 when "01100100010110",
                             7785 when "01100100010111",
                             7783 when "01100100011000",
                             7782 when "01100100011001",
                             7781 when "01100100011010",
                             7780 when "01100100011011",
                             7778 when "01100100011100",
                             7777 when "01100100011101",
                             7776 when "01100100011110",
                             7775 when "01100100011111",
                             7774 when "01100100100000",
                             7772 when "01100100100001",
                             7771 when "01100100100010",
                             7770 when "01100100100011",
                             7769 when "01100100100100",
                             7768 when "01100100100101",
                             7766 when "01100100100110",
                             7765 when "01100100100111",
                             7764 when "01100100101000",
                             7763 when "01100100101001",
                             7762 when "01100100101010",
                             7760 when "01100100101011",
                             7759 when "01100100101100",
                             7758 when "01100100101101",
                             7757 when "01100100101110",
                             7756 when "01100100101111",
                             7754 when "01100100110000",
                             7753 when "01100100110001",
                             7752 when "01100100110010",
                             7751 when "01100100110011",
                             7750 when "01100100110100",
                             7748 when "01100100110101",
                             7747 when "01100100110110",
                             7746 when "01100100110111",
                             7745 when "01100100111000",
                             7744 when "01100100111001",
                             7742 when "01100100111010",
                             7741 when "01100100111011",
                             7740 when "01100100111100",
                             7739 when "01100100111101",
                             7738 when "01100100111110",
                             7736 when "01100100111111",
                             7735 when "01100101000000",
                             7734 when "01100101000001",
                             7733 when "01100101000010",
                             7732 when "01100101000011",
                             7730 when "01100101000100",
                             7729 when "01100101000101",
                             7728 when "01100101000110",
                             7727 when "01100101000111",
                             7726 when "01100101001000",
                             7724 when "01100101001001",
                             7723 when "01100101001010",
                             7722 when "01100101001011",
                             7721 when "01100101001100",
                             7720 when "01100101001101",
                             7718 when "01100101001110",
                             7717 when "01100101001111",
                             7716 when "01100101010000",
                             7715 when "01100101010001",
                             7714 when "01100101010010",
                             7712 when "01100101010011",
                             7711 when "01100101010100",
                             7710 when "01100101010101",
                             7709 when "01100101010110",
                             7708 when "01100101010111",
                             7707 when "01100101011000",
                             7705 when "01100101011001",
                             7704 when "01100101011010",
                             7703 when "01100101011011",
                             7702 when "01100101011100",
                             7701 when "01100101011101",
                             7699 when "01100101011110",
                             7698 when "01100101011111",
                             7697 when "01100101100000",
                             7696 when "01100101100001",
                             7695 when "01100101100010",
                             7693 when "01100101100011",
                             7692 when "01100101100100",
                             7691 when "01100101100101",
                             7690 when "01100101100110",
                             7689 when "01100101100111",
                             7688 when "01100101101000",
                             7686 when "01100101101001",
                             7685 when "01100101101010",
                             7684 when "01100101101011",
                             7683 when "01100101101100",
                             7682 when "01100101101101",
                             7680 when "01100101101110",
                             7679 when "01100101101111",
                             7678 when "01100101110000",
                             7677 when "01100101110001",
                             7676 when "01100101110010",
                             7675 when "01100101110011",
                             7673 when "01100101110100",
                             7672 when "01100101110101",
                             7671 when "01100101110110",
                             7670 when "01100101110111",
                             7669 when "01100101111000",
                             7668 when "01100101111001",
                             7666 when "01100101111010",
                             7665 when "01100101111011",
                             7664 when "01100101111100",
                             7663 when "01100101111101",
                             7662 when "01100101111110",
                             7660 when "01100101111111",
                             7659 when "01100110000000",
                             7658 when "01100110000001",
                             7657 when "01100110000010",
                             7656 when "01100110000011",
                             7655 when "01100110000100",
                             7653 when "01100110000101",
                             7652 when "01100110000110",
                             7651 when "01100110000111",
                             7650 when "01100110001000",
                             7649 when "01100110001001",
                             7648 when "01100110001010",
                             7646 when "01100110001011",
                             7645 when "01100110001100",
                             7644 when "01100110001101",
                             7643 when "01100110001110",
                             7642 when "01100110001111",
                             7641 when "01100110010000",
                             7639 when "01100110010001",
                             7638 when "01100110010010",
                             7637 when "01100110010011",
                             7636 when "01100110010100",
                             7635 when "01100110010101",
                             7634 when "01100110010110",
                             7632 when "01100110010111",
                             7631 when "01100110011000",
                             7630 when "01100110011001",
                             7629 when "01100110011010",
                             7628 when "01100110011011",
                             7627 when "01100110011100",
                             7625 when "01100110011101",
                             7624 when "01100110011110",
                             7623 when "01100110011111",
                             7622 when "01100110100000",
                             7621 when "01100110100001",
                             7620 when "01100110100010",
                             7618 when "01100110100011",
                             7617 when "01100110100100",
                             7616 when "01100110100101",
                             7615 when "01100110100110",
                             7614 when "01100110100111",
                             7613 when "01100110101000",
                             7612 when "01100110101001",
                             7610 when "01100110101010",
                             7609 when "01100110101011",
                             7608 when "01100110101100",
                             7607 when "01100110101101",
                             7606 when "01100110101110",
                             7605 when "01100110101111",
                             7603 when "01100110110000",
                             7602 when "01100110110001",
                             7601 when "01100110110010",
                             7600 when "01100110110011",
                             7599 when "01100110110100",
                             7598 when "01100110110101",
                             7596 when "01100110110110",
                             7595 when "01100110110111",
                             7594 when "01100110111000",
                             7593 when "01100110111001",
                             7592 when "01100110111010",
                             7591 when "01100110111011",
                             7590 when "01100110111100",
                             7588 when "01100110111101",
                             7587 when "01100110111110",
                             7586 when "01100110111111",
                             7585 when "01100111000000",
                             7584 when "01100111000001",
                             7583 when "01100111000010",
                             7582 when "01100111000011",
                             7580 when "01100111000100",
                             7579 when "01100111000101",
                             7578 when "01100111000110",
                             7577 when "01100111000111",
                             7576 when "01100111001000",
                             7575 when "01100111001001",
                             7573 when "01100111001010",
                             7572 when "01100111001011",
                             7571 when "01100111001100",
                             7570 when "01100111001101",
                             7569 when "01100111001110",
                             7568 when "01100111001111",
                             7567 when "01100111010000",
                             7565 when "01100111010001",
                             7564 when "01100111010010",
                             7563 when "01100111010011",
                             7562 when "01100111010100",
                             7561 when "01100111010101",
                             7560 when "01100111010110",
                             7559 when "01100111010111",
                             7557 when "01100111011000",
                             7556 when "01100111011001",
                             7555 when "01100111011010",
                             7554 when "01100111011011",
                             7553 when "01100111011100",
                             7552 when "01100111011101",
                             7551 when "01100111011110",
                             7549 when "01100111011111",
                             7548 when "01100111100000",
                             7547 when "01100111100001",
                             7546 when "01100111100010",
                             7545 when "01100111100011",
                             7544 when "01100111100100",
                             7543 when "01100111100101",
                             7541 when "01100111100110",
                             7540 when "01100111100111",
                             7539 when "01100111101000",
                             7538 when "01100111101001",
                             7537 when "01100111101010",
                             7536 when "01100111101011",
                             7535 when "01100111101100",
                             7534 when "01100111101101",
                             7532 when "01100111101110",
                             7531 when "01100111101111",
                             7530 when "01100111110000",
                             7529 when "01100111110001",
                             7528 when "01100111110010",
                             7527 when "01100111110011",
                             7526 when "01100111110100",
                             7524 when "01100111110101",
                             7523 when "01100111110110",
                             7522 when "01100111110111",
                             7521 when "01100111111000",
                             7520 when "01100111111001",
                             7519 when "01100111111010",
                             7518 when "01100111111011",
                             7517 when "01100111111100",
                             7515 when "01100111111101",
                             7514 when "01100111111110",
                             7513 when "01100111111111",
                             7512 when "01101000000000",
                             7511 when "01101000000001",
                             7510 when "01101000000010",
                             7509 when "01101000000011",
                             7508 when "01101000000100",
                             7506 when "01101000000101",
                             7505 when "01101000000110",
                             7504 when "01101000000111",
                             7503 when "01101000001000",
                             7502 when "01101000001001",
                             7501 when "01101000001010",
                             7500 when "01101000001011",
                             7499 when "01101000001100",
                             7497 when "01101000001101",
                             7496 when "01101000001110",
                             7495 when "01101000001111",
                             7494 when "01101000010000",
                             7493 when "01101000010001",
                             7492 when "01101000010010",
                             7491 when "01101000010011",
                             7490 when "01101000010100",
                             7488 when "01101000010101",
                             7487 when "01101000010110",
                             7486 when "01101000010111",
                             7485 when "01101000011000",
                             7484 when "01101000011001",
                             7483 when "01101000011010",
                             7482 when "01101000011011",
                             7481 when "01101000011100",
                             7479 when "01101000011101",
                             7478 when "01101000011110",
                             7477 when "01101000011111",
                             7476 when "01101000100000",
                             7475 when "01101000100001",
                             7474 when "01101000100010",
                             7473 when "01101000100011",
                             7472 when "01101000100100",
                             7470 when "01101000100101",
                             7469 when "01101000100110",
                             7468 when "01101000100111",
                             7467 when "01101000101000",
                             7466 when "01101000101001",
                             7465 when "01101000101010",
                             7464 when "01101000101011",
                             7463 when "01101000101100",
                             7462 when "01101000101101",
                             7460 when "01101000101110",
                             7459 when "01101000101111",
                             7458 when "01101000110000",
                             7457 when "01101000110001",
                             7456 when "01101000110010",
                             7455 when "01101000110011",
                             7454 when "01101000110100",
                             7453 when "01101000110101",
                             7452 when "01101000110110",
                             7450 when "01101000110111",
                             7449 when "01101000111000",
                             7448 when "01101000111001",
                             7447 when "01101000111010",
                             7446 when "01101000111011",
                             7445 when "01101000111100",
                             7444 when "01101000111101",
                             7443 when "01101000111110",
                             7442 when "01101000111111",
                             7440 when "01101001000000",
                             7439 when "01101001000001",
                             7438 when "01101001000010",
                             7437 when "01101001000011",
                             7436 when "01101001000100",
                             7435 when "01101001000101",
                             7434 when "01101001000110",
                             7433 when "01101001000111",
                             7432 when "01101001001000",
                             7431 when "01101001001001",
                             7429 when "01101001001010",
                             7428 when "01101001001011",
                             7427 when "01101001001100",
                             7426 when "01101001001101",
                             7425 when "01101001001110",
                             7424 when "01101001001111",
                             7423 when "01101001010000",
                             7422 when "01101001010001",
                             7421 when "01101001010010",
                             7419 when "01101001010011",
                             7418 when "01101001010100",
                             7417 when "01101001010101",
                             7416 when "01101001010110",
                             7415 when "01101001010111",
                             7414 when "01101001011000",
                             7413 when "01101001011001",
                             7412 when "01101001011010",
                             7411 when "01101001011011",
                             7410 when "01101001011100",
                             7409 when "01101001011101",
                             7407 when "01101001011110",
                             7406 when "01101001011111",
                             7405 when "01101001100000",
                             7404 when "01101001100001",
                             7403 when "01101001100010",
                             7402 when "01101001100011",
                             7401 when "01101001100100",
                             7400 when "01101001100101",
                             7399 when "01101001100110",
                             7398 when "01101001100111",
                             7396 when "01101001101000",
                             7395 when "01101001101001",
                             7394 when "01101001101010",
                             7393 when "01101001101011",
                             7392 when "01101001101100",
                             7391 when "01101001101101",
                             7390 when "01101001101110",
                             7389 when "01101001101111",
                             7388 when "01101001110000",
                             7387 when "01101001110001",
                             7386 when "01101001110010",
                             7384 when "01101001110011",
                             7383 when "01101001110100",
                             7382 when "01101001110101",
                             7381 when "01101001110110",
                             7380 when "01101001110111",
                             7379 when "01101001111000",
                             7378 when "01101001111001",
                             7377 when "01101001111010",
                             7376 when "01101001111011",
                             7375 when "01101001111100",
                             7374 when "01101001111101",
                             7372 when "01101001111110",
                             7371 when "01101001111111",
                             7370 when "01101010000000",
                             7369 when "01101010000001",
                             7368 when "01101010000010",
                             7367 when "01101010000011",
                             7366 when "01101010000100",
                             7365 when "01101010000101",
                             7364 when "01101010000110",
                             7363 when "01101010000111",
                             7362 when "01101010001000",
                             7361 when "01101010001001",
                             7359 when "01101010001010",
                             7358 when "01101010001011",
                             7357 when "01101010001100",
                             7356 when "01101010001101",
                             7355 when "01101010001110",
                             7354 when "01101010001111",
                             7353 when "01101010010000",
                             7352 when "01101010010001",
                             7351 when "01101010010010",
                             7350 when "01101010010011",
                             7349 when "01101010010100",
                             7348 when "01101010010101",
                             7346 when "01101010010110",
                             7345 when "01101010010111",
                             7344 when "01101010011000",
                             7343 when "01101010011001",
                             7342 when "01101010011010",
                             7341 when "01101010011011",
                             7340 when "01101010011100",
                             7339 when "01101010011101",
                             7338 when "01101010011110",
                             7337 when "01101010011111",
                             7336 when "01101010100000",
                             7335 when "01101010100001",
                             7334 when "01101010100010",
                             7332 when "01101010100011",
                             7331 when "01101010100100",
                             7330 when "01101010100101",
                             7329 when "01101010100110",
                             7328 when "01101010100111",
                             7327 when "01101010101000",
                             7326 when "01101010101001",
                             7325 when "01101010101010",
                             7324 when "01101010101011",
                             7323 when "01101010101100",
                             7322 when "01101010101101",
                             7321 when "01101010101110",
                             7320 when "01101010101111",
                             7319 when "01101010110000",
                             7317 when "01101010110001",
                             7316 when "01101010110010",
                             7315 when "01101010110011",
                             7314 when "01101010110100",
                             7313 when "01101010110101",
                             7312 when "01101010110110",
                             7311 when "01101010110111",
                             7310 when "01101010111000",
                             7309 when "01101010111001",
                             7308 when "01101010111010",
                             7307 when "01101010111011",
                             7306 when "01101010111100",
                             7305 when "01101010111101",
                             7304 when "01101010111110",
                             7302 when "01101010111111",
                             7301 when "01101011000000",
                             7300 when "01101011000001",
                             7299 when "01101011000010",
                             7298 when "01101011000011",
                             7297 when "01101011000100",
                             7296 when "01101011000101",
                             7295 when "01101011000110",
                             7294 when "01101011000111",
                             7293 when "01101011001000",
                             7292 when "01101011001001",
                             7291 when "01101011001010",
                             7290 when "01101011001011",
                             7289 when "01101011001100",
                             7288 when "01101011001101",
                             7287 when "01101011001110",
                             7285 when "01101011001111",
                             7284 when "01101011010000",
                             7283 when "01101011010001",
                             7282 when "01101011010010",
                             7281 when "01101011010011",
                             7280 when "01101011010100",
                             7279 when "01101011010101",
                             7278 when "01101011010110",
                             7277 when "01101011010111",
                             7276 when "01101011011000",
                             7275 when "01101011011001",
                             7274 when "01101011011010",
                             7273 when "01101011011011",
                             7272 when "01101011011100",
                             7271 when "01101011011101",
                             7270 when "01101011011110",
                             7268 when "01101011011111",
                             7267 when "01101011100000",
                             7266 when "01101011100001",
                             7265 when "01101011100010",
                             7264 when "01101011100011",
                             7263 when "01101011100100",
                             7262 when "01101011100101",
                             7261 when "01101011100110",
                             7260 when "01101011100111",
                             7259 when "01101011101000",
                             7258 when "01101011101001",
                             7257 when "01101011101010",
                             7256 when "01101011101011",
                             7255 when "01101011101100",
                             7254 when "01101011101101",
                             7253 when "01101011101110",
                             7252 when "01101011101111",
                             7251 when "01101011110000",
                             7250 when "01101011110001",
                             7248 when "01101011110010",
                             7247 when "01101011110011",
                             7246 when "01101011110100",
                             7245 when "01101011110101",
                             7244 when "01101011110110",
                             7243 when "01101011110111",
                             7242 when "01101011111000",
                             7241 when "01101011111001",
                             7240 when "01101011111010",
                             7239 when "01101011111011",
                             7238 when "01101011111100",
                             7237 when "01101011111101",
                             7236 when "01101011111110",
                             7235 when "01101011111111",
                             7234 when "01101100000000",
                             7233 when "01101100000001",
                             7232 when "01101100000010",
                             7231 when "01101100000011",
                             7230 when "01101100000100",
                             7229 when "01101100000101",
                             7228 when "01101100000110",
                             7226 when "01101100000111",
                             7225 when "01101100001000",
                             7224 when "01101100001001",
                             7223 when "01101100001010",
                             7222 when "01101100001011",
                             7221 when "01101100001100",
                             7220 when "01101100001101",
                             7219 when "01101100001110",
                             7218 when "01101100001111",
                             7217 when "01101100010000",
                             7216 when "01101100010001",
                             7215 when "01101100010010",
                             7214 when "01101100010011",
                             7213 when "01101100010100",
                             7212 when "01101100010101",
                             7211 when "01101100010110",
                             7210 when "01101100010111",
                             7209 when "01101100011000",
                             7208 when "01101100011001",
                             7207 when "01101100011010",
                             7206 when "01101100011011",
                             7205 when "01101100011100",
                             7204 when "01101100011101",
                             7203 when "01101100011110",
                             7201 when "01101100011111",
                             7200 when "01101100100000",
                             7199 when "01101100100001",
                             7198 when "01101100100010",
                             7197 when "01101100100011",
                             7196 when "01101100100100",
                             7195 when "01101100100101",
                             7194 when "01101100100110",
                             7193 when "01101100100111",
                             7192 when "01101100101000",
                             7191 when "01101100101001",
                             7190 when "01101100101010",
                             7189 when "01101100101011",
                             7188 when "01101100101100",
                             7187 when "01101100101101",
                             7186 when "01101100101110",
                             7185 when "01101100101111",
                             7184 when "01101100110000",
                             7183 when "01101100110001",
                             7182 when "01101100110010",
                             7181 when "01101100110011",
                             7180 when "01101100110100",
                             7179 when "01101100110101",
                             7178 when "01101100110110",
                             7177 when "01101100110111",
                             7176 when "01101100111000",
                             7175 when "01101100111001",
                             7174 when "01101100111010",
                             7173 when "01101100111011",
                             7172 when "01101100111100",
                             7171 when "01101100111101",
                             7169 when "01101100111110",
                             7168 when "01101100111111",
                             7167 when "01101101000000",
                             7166 when "01101101000001",
                             7165 when "01101101000010",
                             7164 when "01101101000011",
                             7163 when "01101101000100",
                             7162 when "01101101000101",
                             7161 when "01101101000110",
                             7160 when "01101101000111",
                             7159 when "01101101001000",
                             7158 when "01101101001001",
                             7157 when "01101101001010",
                             7156 when "01101101001011",
                             7155 when "01101101001100",
                             7154 when "01101101001101",
                             7153 when "01101101001110",
                             7152 when "01101101001111",
                             7151 when "01101101010000",
                             7150 when "01101101010001",
                             7149 when "01101101010010",
                             7148 when "01101101010011",
                             7147 when "01101101010100",
                             7146 when "01101101010101",
                             7145 when "01101101010110",
                             7144 when "01101101010111",
                             7143 when "01101101011000",
                             7142 when "01101101011001",
                             7141 when "01101101011010",
                             7140 when "01101101011011",
                             7139 when "01101101011100",
                             7138 when "01101101011101",
                             7137 when "01101101011110",
                             7136 when "01101101011111",
                             7135 when "01101101100000",
                             7134 when "01101101100001",
                             7133 when "01101101100010",
                             7132 when "01101101100011",
                             7131 when "01101101100100",
                             7130 when "01101101100101",
                             7129 when "01101101100110",
                             7128 when "01101101100111",
                             7127 when "01101101101000",
                             7126 when "01101101101001",
                             7125 when "01101101101010",
                             7124 when "01101101101011",
                             7123 when "01101101101100",
                             7121 when "01101101101101",
                             7120 when "01101101101110",
                             7119 when "01101101101111",
                             7118 when "01101101110000",
                             7117 when "01101101110001",
                             7116 when "01101101110010",
                             7115 when "01101101110011",
                             7114 when "01101101110100",
                             7113 when "01101101110101",
                             7112 when "01101101110110",
                             7111 when "01101101110111",
                             7110 when "01101101111000",
                             7109 when "01101101111001",
                             7108 when "01101101111010",
                             7107 when "01101101111011",
                             7106 when "01101101111100",
                             7105 when "01101101111101",
                             7104 when "01101101111110",
                             7103 when "01101101111111",
                             7102 when "01101110000000",
                             7101 when "01101110000001",
                             7100 when "01101110000010",
                             7099 when "01101110000011",
                             7098 when "01101110000100",
                             7097 when "01101110000101",
                             7096 when "01101110000110",
                             7095 when "01101110000111",
                             7094 when "01101110001000",
                             7093 when "01101110001001",
                             7092 when "01101110001010",
                             7091 when "01101110001011",
                             7090 when "01101110001100",
                             7089 when "01101110001101",
                             7088 when "01101110001110",
                             7087 when "01101110001111",
                             7086 when "01101110010000",
                             7085 when "01101110010001",
                             7084 when "01101110010010",
                             7083 when "01101110010011",
                             7082 when "01101110010100",
                             7081 when "01101110010101",
                             7080 when "01101110010110",
                             7079 when "01101110010111",
                             7078 when "01101110011000",
                             7077 when "01101110011001",
                             7076 when "01101110011010",
                             7075 when "01101110011011",
                             7074 when "01101110011100",
                             7073 when "01101110011101",
                             7072 when "01101110011110",
                             7071 when "01101110011111",
                             7070 when "01101110100000",
                             7069 when "01101110100001",
                             7068 when "01101110100010",
                             7067 when "01101110100011",
                             7066 when "01101110100100",
                             7065 when "01101110100101",
                             7064 when "01101110100110",
                             7063 when "01101110100111",
                             7062 when "01101110101000",
                             7061 when "01101110101001",
                             7060 when "01101110101010",
                             7059 when "01101110101011",
                             7058 when "01101110101100",
                             7057 when "01101110101101",
                             7056 when "01101110101110",
                             7055 when "01101110101111",
                             7054 when "01101110110000",
                             7053 when "01101110110001",
                             7052 when "01101110110010",
                             7051 when "01101110110011",
                             7050 when "01101110110100",
                             7049 when "01101110110101",
                             7048 when "01101110110110",
                             7047 when "01101110110111",
                             7046 when "01101110111000",
                             7045 when "01101110111001",
                             7044 when "01101110111010",
                             7043 when "01101110111011",
                             7042 when "01101110111100",
                             7041 when "01101110111101",
                             7040 when "01101110111110",
                             7039 when "01101110111111",
                             7038 when "01101111000000",
                             7037 when "01101111000001",
                             7036 when "01101111000010",
                             7035 when "01101111000011",
                             7034 when "01101111000100",
                             7033 when "01101111000101",
                             7032 when "01101111000110",
                             7031 when "01101111000111",
                             7030 when "01101111001000",
                             7029 when "01101111001001",
                             7028 when "01101111001010",
                             7027 when "01101111001011",
                             7026 when "01101111001100",
                             7025 when "01101111001101",
                             7024 when "01101111001110",
                             7023 when "01101111001111",
                             7022 when "01101111010000",
                             7021 when "01101111010001",
                             7020 when "01101111010010",
                             7020 when "01101111010011",
                             7019 when "01101111010100",
                             7018 when "01101111010101",
                             7017 when "01101111010110",
                             7016 when "01101111010111",
                             7015 when "01101111011000",
                             7014 when "01101111011001",
                             7013 when "01101111011010",
                             7012 when "01101111011011",
                             7011 when "01101111011100",
                             7010 when "01101111011101",
                             7009 when "01101111011110",
                             7008 when "01101111011111",
                             7007 when "01101111100000",
                             7006 when "01101111100001",
                             7005 when "01101111100010",
                             7004 when "01101111100011",
                             7003 when "01101111100100",
                             7002 when "01101111100101",
                             7001 when "01101111100110",
                             7000 when "01101111100111",
                             6999 when "01101111101000",
                             6998 when "01101111101001",
                             6997 when "01101111101010",
                             6996 when "01101111101011",
                             6995 when "01101111101100",
                             6994 when "01101111101101",
                             6993 when "01101111101110",
                             6992 when "01101111101111",
                             6991 when "01101111110000",
                             6990 when "01101111110001",
                             6989 when "01101111110010",
                             6988 when "01101111110011",
                             6987 when "01101111110100",
                             6986 when "01101111110101",
                             6985 when "01101111110110",
                             6984 when "01101111110111",
                             6983 when "01101111111000",
                             6982 when "01101111111001",
                             6981 when "01101111111010",
                             6980 when "01101111111011",
                             6979 when "01101111111100",
                             6978 when "01101111111101",
                             6977 when "01101111111110",
                             6976 when "01101111111111",
                             6975 when "01110000000000",
                             6974 when "01110000000001",
                             6974 when "01110000000010",
                             6973 when "01110000000011",
                             6972 when "01110000000100",
                             6971 when "01110000000101",
                             6970 when "01110000000110",
                             6969 when "01110000000111",
                             6968 when "01110000001000",
                             6967 when "01110000001001",
                             6966 when "01110000001010",
                             6965 when "01110000001011",
                             6964 when "01110000001100",
                             6963 when "01110000001101",
                             6962 when "01110000001110",
                             6961 when "01110000001111",
                             6960 when "01110000010000",
                             6959 when "01110000010001",
                             6958 when "01110000010010",
                             6957 when "01110000010011",
                             6956 when "01110000010100",
                             6955 when "01110000010101",
                             6954 when "01110000010110",
                             6953 when "01110000010111",
                             6952 when "01110000011000",
                             6951 when "01110000011001",
                             6950 when "01110000011010",
                             6949 when "01110000011011",
                             6948 when "01110000011100",
                             6947 when "01110000011101",
                             6946 when "01110000011110",
                             6945 when "01110000011111",
                             6944 when "01110000100000",
                             6943 when "01110000100001",
                             6943 when "01110000100010",
                             6942 when "01110000100011",
                             6941 when "01110000100100",
                             6940 when "01110000100101",
                             6939 when "01110000100110",
                             6938 when "01110000100111",
                             6937 when "01110000101000",
                             6936 when "01110000101001",
                             6935 when "01110000101010",
                             6934 when "01110000101011",
                             6933 when "01110000101100",
                             6932 when "01110000101101",
                             6931 when "01110000101110",
                             6930 when "01110000101111",
                             6929 when "01110000110000",
                             6928 when "01110000110001",
                             6927 when "01110000110010",
                             6926 when "01110000110011",
                             6925 when "01110000110100",
                             6924 when "01110000110101",
                             6923 when "01110000110110",
                             6922 when "01110000110111",
                             6921 when "01110000111000",
                             6920 when "01110000111001",
                             6919 when "01110000111010",
                             6919 when "01110000111011",
                             6918 when "01110000111100",
                             6917 when "01110000111101",
                             6916 when "01110000111110",
                             6915 when "01110000111111",
                             6914 when "01110001000000",
                             6913 when "01110001000001",
                             6912 when "01110001000010",
                             6911 when "01110001000011",
                             6910 when "01110001000100",
                             6909 when "01110001000101",
                             6908 when "01110001000110",
                             6907 when "01110001000111",
                             6906 when "01110001001000",
                             6905 when "01110001001001",
                             6904 when "01110001001010",
                             6903 when "01110001001011",
                             6902 when "01110001001100",
                             6901 when "01110001001101",
                             6900 when "01110001001110",
                             6899 when "01110001001111",
                             6898 when "01110001010000",
                             6898 when "01110001010001",
                             6897 when "01110001010010",
                             6896 when "01110001010011",
                             6895 when "01110001010100",
                             6894 when "01110001010101",
                             6893 when "01110001010110",
                             6892 when "01110001010111",
                             6891 when "01110001011000",
                             6890 when "01110001011001",
                             6889 when "01110001011010",
                             6888 when "01110001011011",
                             6887 when "01110001011100",
                             6886 when "01110001011101",
                             6885 when "01110001011110",
                             6884 when "01110001011111",
                             6883 when "01110001100000",
                             6882 when "01110001100001",
                             6881 when "01110001100010",
                             6880 when "01110001100011",
                             6879 when "01110001100100",
                             6879 when "01110001100101",
                             6878 when "01110001100110",
                             6877 when "01110001100111",
                             6876 when "01110001101000",
                             6875 when "01110001101001",
                             6874 when "01110001101010",
                             6873 when "01110001101011",
                             6872 when "01110001101100",
                             6871 when "01110001101101",
                             6870 when "01110001101110",
                             6869 when "01110001101111",
                             6868 when "01110001110000",
                             6867 when "01110001110001",
                             6866 when "01110001110010",
                             6865 when "01110001110011",
                             6864 when "01110001110100",
                             6863 when "01110001110101",
                             6862 when "01110001110110",
                             6862 when "01110001110111",
                             6861 when "01110001111000",
                             6860 when "01110001111001",
                             6859 when "01110001111010",
                             6858 when "01110001111011",
                             6857 when "01110001111100",
                             6856 when "01110001111101",
                             6855 when "01110001111110",
                             6854 when "01110001111111",
                             6853 when "01110010000000",
                             6852 when "01110010000001",
                             6851 when "01110010000010",
                             6850 when "01110010000011",
                             6849 when "01110010000100",
                             6848 when "01110010000101",
                             6847 when "01110010000110",
                             6847 when "01110010000111",
                             6846 when "01110010001000",
                             6845 when "01110010001001",
                             6844 when "01110010001010",
                             6843 when "01110010001011",
                             6842 when "01110010001100",
                             6841 when "01110010001101",
                             6840 when "01110010001110",
                             6839 when "01110010001111",
                             6838 when "01110010010000",
                             6837 when "01110010010001",
                             6836 when "01110010010010",
                             6835 when "01110010010011",
                             6834 when "01110010010100",
                             6833 when "01110010010101",
                             6832 when "01110010010110",
                             6832 when "01110010010111",
                             6831 when "01110010011000",
                             6830 when "01110010011001",
                             6829 when "01110010011010",
                             6828 when "01110010011011",
                             6827 when "01110010011100",
                             6826 when "01110010011101",
                             6825 when "01110010011110",
                             6824 when "01110010011111",
                             6823 when "01110010100000",
                             6822 when "01110010100001",
                             6821 when "01110010100010",
                             6820 when "01110010100011",
                             6819 when "01110010100100",
                             6818 when "01110010100101",
                             6818 when "01110010100110",
                             6817 when "01110010100111",
                             6816 when "01110010101000",
                             6815 when "01110010101001",
                             6814 when "01110010101010",
                             6813 when "01110010101011",
                             6812 when "01110010101100",
                             6811 when "01110010101101",
                             6810 when "01110010101110",
                             6809 when "01110010101111",
                             6808 when "01110010110000",
                             6807 when "01110010110001",
                             6806 when "01110010110010",
                             6805 when "01110010110011",
                             6805 when "01110010110100",
                             6804 when "01110010110101",
                             6803 when "01110010110110",
                             6802 when "01110010110111",
                             6801 when "01110010111000",
                             6800 when "01110010111001",
                             6799 when "01110010111010",
                             6798 when "01110010111011",
                             6797 when "01110010111100",
                             6796 when "01110010111101",
                             6795 when "01110010111110",
                             6794 when "01110010111111",
                             6793 when "01110011000000",
                             6793 when "01110011000001",
                             6792 when "01110011000010",
                             6791 when "01110011000011",
                             6790 when "01110011000100",
                             6789 when "01110011000101",
                             6788 when "01110011000110",
                             6787 when "01110011000111",
                             6786 when "01110011001000",
                             6785 when "01110011001001",
                             6784 when "01110011001010",
                             6783 when "01110011001011",
                             6782 when "01110011001100",
                             6782 when "01110011001101",
                             6781 when "01110011001110",
                             6780 when "01110011001111",
                             6779 when "01110011010000",
                             6778 when "01110011010001",
                             6777 when "01110011010010",
                             6776 when "01110011010011",
                             6775 when "01110011010100",
                             6774 when "01110011010101",
                             6773 when "01110011010110",
                             6772 when "01110011010111",
                             6771 when "01110011011000",
                             6770 when "01110011011001",
                             6770 when "01110011011010",
                             6769 when "01110011011011",
                             6768 when "01110011011100",
                             6767 when "01110011011101",
                             6766 when "01110011011110",
                             6765 when "01110011011111",
                             6764 when "01110011100000",
                             6763 when "01110011100001",
                             6762 when "01110011100010",
                             6761 when "01110011100011",
                             6760 when "01110011100100",
                             6759 when "01110011100101",
                             6759 when "01110011100110",
                             6758 when "01110011100111",
                             6757 when "01110011101000",
                             6756 when "01110011101001",
                             6755 when "01110011101010",
                             6754 when "01110011101011",
                             6753 when "01110011101100",
                             6752 when "01110011101101",
                             6751 when "01110011101110",
                             6750 when "01110011101111",
                             6749 when "01110011110000",
                             6749 when "01110011110001",
                             6748 when "01110011110010",
                             6747 when "01110011110011",
                             6746 when "01110011110100",
                             6745 when "01110011110101",
                             6744 when "01110011110110",
                             6743 when "01110011110111",
                             6742 when "01110011111000",
                             6741 when "01110011111001",
                             6740 when "01110011111010",
                             6739 when "01110011111011",
                             6739 when "01110011111100",
                             6738 when "01110011111101",
                             6737 when "01110011111110",
                             6736 when "01110011111111",
                             6735 when "01110100000000",
                             6734 when "01110100000001",
                             6733 when "01110100000010",
                             6732 when "01110100000011",
                             6731 when "01110100000100",
                             6730 when "01110100000101",
                             6729 when "01110100000110",
                             6729 when "01110100000111",
                             6728 when "01110100001000",
                             6727 when "01110100001001",
                             6726 when "01110100001010",
                             6725 when "01110100001011",
                             6724 when "01110100001100",
                             6723 when "01110100001101",
                             6722 when "01110100001110",
                             6721 when "01110100001111",
                             6720 when "01110100010000",
                             6720 when "01110100010001",
                             6719 when "01110100010010",
                             6718 when "01110100010011",
                             6717 when "01110100010100",
                             6716 when "01110100010101",
                             6715 when "01110100010110",
                             6714 when "01110100010111",
                             6713 when "01110100011000",
                             6712 when "01110100011001",
                             6711 when "01110100011010",
                             6711 when "01110100011011",
                             6710 when "01110100011100",
                             6709 when "01110100011101",
                             6708 when "01110100011110",
                             6707 when "01110100011111",
                             6706 when "01110100100000",
                             6705 when "01110100100001",
                             6704 when "01110100100010",
                             6703 when "01110100100011",
                             6702 when "01110100100100",
                             6702 when "01110100100101",
                             6701 when "01110100100110",
                             6700 when "01110100100111",
                             6699 when "01110100101000",
                             6698 when "01110100101001",
                             6697 when "01110100101010",
                             6696 when "01110100101011",
                             6695 when "01110100101100",
                             6694 when "01110100101101",
                             6693 when "01110100101110",
                             6693 when "01110100101111",
                             6692 when "01110100110000",
                             6691 when "01110100110001",
                             6690 when "01110100110010",
                             6689 when "01110100110011",
                             6688 when "01110100110100",
                             6687 when "01110100110101",
                             6686 when "01110100110110",
                             6685 when "01110100110111",
                             6684 when "01110100111000",
                             6684 when "01110100111001",
                             6683 when "01110100111010",
                             6682 when "01110100111011",
                             6681 when "01110100111100",
                             6680 when "01110100111101",
                             6679 when "01110100111110",
                             6678 when "01110100111111",
                             6677 when "01110101000000",
                             6676 when "01110101000001",
                             6676 when "01110101000010",
                             6675 when "01110101000011",
                             6674 when "01110101000100",
                             6673 when "01110101000101",
                             6672 when "01110101000110",
                             6671 when "01110101000111",
                             6670 when "01110101001000",
                             6669 when "01110101001001",
                             6668 when "01110101001010",
                             6668 when "01110101001011",
                             6667 when "01110101001100",
                             6666 when "01110101001101",
                             6665 when "01110101001110",
                             6664 when "01110101001111",
                             6663 when "01110101010000",
                             6662 when "01110101010001",
                             6661 when "01110101010010",
                             6660 when "01110101010011",
                             6660 when "01110101010100",
                             6659 when "01110101010101",
                             6658 when "01110101010110",
                             6657 when "01110101010111",
                             6656 when "01110101011000",
                             6655 when "01110101011001",
                             6654 when "01110101011010",
                             6653 when "01110101011011",
                             6652 when "01110101011100",
                             6652 when "01110101011101",
                             6651 when "01110101011110",
                             6650 when "01110101011111",
                             6649 when "01110101100000",
                             6648 when "01110101100001",
                             6647 when "01110101100010",
                             6646 when "01110101100011",
                             6645 when "01110101100100",
                             6645 when "01110101100101",
                             6644 when "01110101100110",
                             6643 when "01110101100111",
                             6642 when "01110101101000",
                             6641 when "01110101101001",
                             6640 when "01110101101010",
                             6639 when "01110101101011",
                             6638 when "01110101101100",
                             6637 when "01110101101101",
                             6637 when "01110101101110",
                             6636 when "01110101101111",
                             6635 when "01110101110000",
                             6634 when "01110101110001",
                             6633 when "01110101110010",
                             6632 when "01110101110011",
                             6631 when "01110101110100",
                             6630 when "01110101110101",
                             6630 when "01110101110110",
                             6629 when "01110101110111",
                             6628 when "01110101111000",
                             6627 when "01110101111001",
                             6626 when "01110101111010",
                             6625 when "01110101111011",
                             6624 when "01110101111100",
                             6623 when "01110101111101",
                             6623 when "01110101111110",
                             6622 when "01110101111111",
                             6621 when "01110110000000",
                             6620 when "01110110000001",
                             6619 when "01110110000010",
                             6618 when "01110110000011",
                             6617 when "01110110000100",
                             6616 when "01110110000101",
                             6616 when "01110110000110",
                             6615 when "01110110000111",
                             6614 when "01110110001000",
                             6613 when "01110110001001",
                             6612 when "01110110001010",
                             6611 when "01110110001011",
                             6610 when "01110110001100",
                             6609 when "01110110001101",
                             6609 when "01110110001110",
                             6608 when "01110110001111",
                             6607 when "01110110010000",
                             6606 when "01110110010001",
                             6605 when "01110110010010",
                             6604 when "01110110010011",
                             6603 when "01110110010100",
                             6602 when "01110110010101",
                             6602 when "01110110010110",
                             6601 when "01110110010111",
                             6600 when "01110110011000",
                             6599 when "01110110011001",
                             6598 when "01110110011010",
                             6597 when "01110110011011",
                             6596 when "01110110011100",
                             6595 when "01110110011101",
                             6595 when "01110110011110",
                             6594 when "01110110011111",
                             6593 when "01110110100000",
                             6592 when "01110110100001",
                             6591 when "01110110100010",
                             6590 when "01110110100011",
                             6589 when "01110110100100",
                             6588 when "01110110100101",
                             6588 when "01110110100110",
                             6587 when "01110110100111",
                             6586 when "01110110101000",
                             6585 when "01110110101001",
                             6584 when "01110110101010",
                             6583 when "01110110101011",
                             6582 when "01110110101100",
                             6582 when "01110110101101",
                             6581 when "01110110101110",
                             6580 when "01110110101111",
                             6579 when "01110110110000",
                             6578 when "01110110110001",
                             6577 when "01110110110010",
                             6576 when "01110110110011",
                             6575 when "01110110110100",
                             6575 when "01110110110101",
                             6574 when "01110110110110",
                             6573 when "01110110110111",
                             6572 when "01110110111000",
                             6571 when "01110110111001",
                             6570 when "01110110111010",
                             6569 when "01110110111011",
                             6569 when "01110110111100",
                             6568 when "01110110111101",
                             6567 when "01110110111110",
                             6566 when "01110110111111",
                             6565 when "01110111000000",
                             6564 when "01110111000001",
                             6563 when "01110111000010",
                             6563 when "01110111000011",
                             6562 when "01110111000100",
                             6561 when "01110111000101",
                             6560 when "01110111000110",
                             6559 when "01110111000111",
                             6558 when "01110111001000",
                             6557 when "01110111001001",
                             6557 when "01110111001010",
                             6556 when "01110111001011",
                             6555 when "01110111001100",
                             6554 when "01110111001101",
                             6553 when "01110111001110",
                             6552 when "01110111001111",
                             6551 when "01110111010000",
                             6551 when "01110111010001",
                             6550 when "01110111010010",
                             6549 when "01110111010011",
                             6548 when "01110111010100",
                             6547 when "01110111010101",
                             6546 when "01110111010110",
                             6545 when "01110111010111",
                             6545 when "01110111011000",
                             6544 when "01110111011001",
                             6543 when "01110111011010",
                             6542 when "01110111011011",
                             6541 when "01110111011100",
                             6540 when "01110111011101",
                             6539 when "01110111011110",
                             6539 when "01110111011111",
                             6538 when "01110111100000",
                             6537 when "01110111100001",
                             6536 when "01110111100010",
                             6535 when "01110111100011",
                             6534 when "01110111100100",
                             6533 when "01110111100101",
                             6533 when "01110111100110",
                             6532 when "01110111100111",
                             6531 when "01110111101000",
                             6530 when "01110111101001",
                             6529 when "01110111101010",
                             6528 when "01110111101011",
                             6527 when "01110111101100",
                             6527 when "01110111101101",
                             6526 when "01110111101110",
                             6525 when "01110111101111",
                             6524 when "01110111110000",
                             6523 when "01110111110001",
                             6522 when "01110111110010",
                             6521 when "01110111110011",
                             6521 when "01110111110100",
                             6520 when "01110111110101",
                             6519 when "01110111110110",
                             6518 when "01110111110111",
                             6517 when "01110111111000",
                             6516 when "01110111111001",
                             6516 when "01110111111010",
                             6515 when "01110111111011",
                             6514 when "01110111111100",
                             6513 when "01110111111101",
                             6512 when "01110111111110",
                             6511 when "01110111111111",
                             6510 when "01111000000000",
                             6510 when "01111000000001",
                             6509 when "01111000000010",
                             6508 when "01111000000011",
                             6507 when "01111000000100",
                             6506 when "01111000000101",
                             6505 when "01111000000110",
                             6504 when "01111000000111",
                             6504 when "01111000001000",
                             6503 when "01111000001001",
                             6502 when "01111000001010",
                             6501 when "01111000001011",
                             6500 when "01111000001100",
                             6499 when "01111000001101",
                             6499 when "01111000001110",
                             6498 when "01111000001111",
                             6497 when "01111000010000",
                             6496 when "01111000010001",
                             6495 when "01111000010010",
                             6494 when "01111000010011",
                             6494 when "01111000010100",
                             6493 when "01111000010101",
                             6492 when "01111000010110",
                             6491 when "01111000010111",
                             6490 when "01111000011000",
                             6489 when "01111000011001",
                             6488 when "01111000011010",
                             6488 when "01111000011011",
                             6487 when "01111000011100",
                             6486 when "01111000011101",
                             6485 when "01111000011110",
                             6484 when "01111000011111",
                             6483 when "01111000100000",
                             6483 when "01111000100001",
                             6482 when "01111000100010",
                             6481 when "01111000100011",
                             6480 when "01111000100100",
                             6479 when "01111000100101",
                             6478 when "01111000100110",
                             6478 when "01111000100111",
                             6477 when "01111000101000",
                             6476 when "01111000101001",
                             6475 when "01111000101010",
                             6474 when "01111000101011",
                             6473 when "01111000101100",
                             6472 when "01111000101101",
                             6472 when "01111000101110",
                             6471 when "01111000101111",
                             6470 when "01111000110000",
                             6469 when "01111000110001",
                             6468 when "01111000110010",
                             6467 when "01111000110011",
                             6467 when "01111000110100",
                             6466 when "01111000110101",
                             6465 when "01111000110110",
                             6464 when "01111000110111",
                             6463 when "01111000111000",
                             6462 when "01111000111001",
                             6462 when "01111000111010",
                             6461 when "01111000111011",
                             6460 when "01111000111100",
                             6459 when "01111000111101",
                             6458 when "01111000111110",
                             6457 when "01111000111111",
                             6457 when "01111001000000",
                             6456 when "01111001000001",
                             6455 when "01111001000010",
                             6454 when "01111001000011",
                             6453 when "01111001000100",
                             6452 when "01111001000101",
                             6452 when "01111001000110",
                             6451 when "01111001000111",
                             6450 when "01111001001000",
                             6449 when "01111001001001",
                             6448 when "01111001001010",
                             6447 when "01111001001011",
                             6447 when "01111001001100",
                             6446 when "01111001001101",
                             6445 when "01111001001110",
                             6444 when "01111001001111",
                             6443 when "01111001010000",
                             6442 when "01111001010001",
                             6442 when "01111001010010",
                             6441 when "01111001010011",
                             6440 when "01111001010100",
                             6439 when "01111001010101",
                             6438 when "01111001010110",
                             6437 when "01111001010111",
                             6437 when "01111001011000",
                             6436 when "01111001011001",
                             6435 when "01111001011010",
                             6434 when "01111001011011",
                             6433 when "01111001011100",
                             6433 when "01111001011101",
                             6432 when "01111001011110",
                             6431 when "01111001011111",
                             6430 when "01111001100000",
                             6429 when "01111001100001",
                             6428 when "01111001100010",
                             6428 when "01111001100011",
                             6427 when "01111001100100",
                             6426 when "01111001100101",
                             6425 when "01111001100110",
                             6424 when "01111001100111",
                             6423 when "01111001101000",
                             6423 when "01111001101001",
                             6422 when "01111001101010",
                             6421 when "01111001101011",
                             6420 when "01111001101100",
                             6419 when "01111001101101",
                             6418 when "01111001101110",
                             6418 when "01111001101111",
                             6417 when "01111001110000",
                             6416 when "01111001110001",
                             6415 when "01111001110010",
                             6414 when "01111001110011",
                             6414 when "01111001110100",
                             6413 when "01111001110101",
                             6412 when "01111001110110",
                             6411 when "01111001110111",
                             6410 when "01111001111000",
                             6409 when "01111001111001",
                             6409 when "01111001111010",
                             6408 when "01111001111011",
                             6407 when "01111001111100",
                             6406 when "01111001111101",
                             6405 when "01111001111110",
                             6405 when "01111001111111",
                             6404 when "01111010000000",
                             6403 when "01111010000001",
                             6402 when "01111010000010",
                             6401 when "01111010000011",
                             6400 when "01111010000100",
                             6400 when "01111010000101",
                             6399 when "01111010000110",
                             6398 when "01111010000111",
                             6397 when "01111010001000",
                             6396 when "01111010001001",
                             6395 when "01111010001010",
                             6395 when "01111010001011",
                             6394 when "01111010001100",
                             6393 when "01111010001101",
                             6392 when "01111010001110",
                             6391 when "01111010001111",
                             6391 when "01111010010000",
                             6390 when "01111010010001",
                             6389 when "01111010010010",
                             6388 when "01111010010011",
                             6387 when "01111010010100",
                             6387 when "01111010010101",
                             6386 when "01111010010110",
                             6385 when "01111010010111",
                             6384 when "01111010011000",
                             6383 when "01111010011001",
                             6382 when "01111010011010",
                             6382 when "01111010011011",
                             6381 when "01111010011100",
                             6380 when "01111010011101",
                             6379 when "01111010011110",
                             6378 when "01111010011111",
                             6378 when "01111010100000",
                             6377 when "01111010100001",
                             6376 when "01111010100010",
                             6375 when "01111010100011",
                             6374 when "01111010100100",
                             6373 when "01111010100101",
                             6373 when "01111010100110",
                             6372 when "01111010100111",
                             6371 when "01111010101000",
                             6370 when "01111010101001",
                             6369 when "01111010101010",
                             6369 when "01111010101011",
                             6368 when "01111010101100",
                             6367 when "01111010101101",
                             6366 when "01111010101110",
                             6365 when "01111010101111",
                             6365 when "01111010110000",
                             6364 when "01111010110001",
                             6363 when "01111010110010",
                             6362 when "01111010110011",
                             6361 when "01111010110100",
                             6361 when "01111010110101",
                             6360 when "01111010110110",
                             6359 when "01111010110111",
                             6358 when "01111010111000",
                             6357 when "01111010111001",
                             6356 when "01111010111010",
                             6356 when "01111010111011",
                             6355 when "01111010111100",
                             6354 when "01111010111101",
                             6353 when "01111010111110",
                             6352 when "01111010111111",
                             6352 when "01111011000000",
                             6351 when "01111011000001",
                             6350 when "01111011000010",
                             6349 when "01111011000011",
                             6348 when "01111011000100",
                             6348 when "01111011000101",
                             6347 when "01111011000110",
                             6346 when "01111011000111",
                             6345 when "01111011001000",
                             6344 when "01111011001001",
                             6344 when "01111011001010",
                             6343 when "01111011001011",
                             6342 when "01111011001100",
                             6341 when "01111011001101",
                             6340 when "01111011001110",
                             6340 when "01111011001111",
                             6339 when "01111011010000",
                             6338 when "01111011010001",
                             6337 when "01111011010010",
                             6336 when "01111011010011",
                             6336 when "01111011010100",
                             6335 when "01111011010101",
                             6334 when "01111011010110",
                             6333 when "01111011010111",
                             6332 when "01111011011000",
                             6332 when "01111011011001",
                             6331 when "01111011011010",
                             6330 when "01111011011011",
                             6329 when "01111011011100",
                             6328 when "01111011011101",
                             6328 when "01111011011110",
                             6327 when "01111011011111",
                             6326 when "01111011100000",
                             6325 when "01111011100001",
                             6324 when "01111011100010",
                             6324 when "01111011100011",
                             6323 when "01111011100100",
                             6322 when "01111011100101",
                             6321 when "01111011100110",
                             6320 when "01111011100111",
                             6320 when "01111011101000",
                             6319 when "01111011101001",
                             6318 when "01111011101010",
                             6317 when "01111011101011",
                             6316 when "01111011101100",
                             6316 when "01111011101101",
                             6315 when "01111011101110",
                             6314 when "01111011101111",
                             6313 when "01111011110000",
                             6312 when "01111011110001",
                             6312 when "01111011110010",
                             6311 when "01111011110011",
                             6310 when "01111011110100",
                             6309 when "01111011110101",
                             6308 when "01111011110110",
                             6308 when "01111011110111",
                             6307 when "01111011111000",
                             6306 when "01111011111001",
                             6305 when "01111011111010",
                             6304 when "01111011111011",
                             6304 when "01111011111100",
                             6303 when "01111011111101",
                             6302 when "01111011111110",
                             6301 when "01111011111111",
                             6300 when "01111100000000",
                             6300 when "01111100000001",
                             6299 when "01111100000010",
                             6298 when "01111100000011",
                             6297 when "01111100000100",
                             6296 when "01111100000101",
                             6296 when "01111100000110",
                             6295 when "01111100000111",
                             6294 when "01111100001000",
                             6293 when "01111100001001",
                             6292 when "01111100001010",
                             6292 when "01111100001011",
                             6291 when "01111100001100",
                             6290 when "01111100001101",
                             6289 when "01111100001110",
                             6289 when "01111100001111",
                             6288 when "01111100010000",
                             6287 when "01111100010001",
                             6286 when "01111100010010",
                             6285 when "01111100010011",
                             6285 when "01111100010100",
                             6284 when "01111100010101",
                             6283 when "01111100010110",
                             6282 when "01111100010111",
                             6281 when "01111100011000",
                             6281 when "01111100011001",
                             6280 when "01111100011010",
                             6279 when "01111100011011",
                             6278 when "01111100011100",
                             6277 when "01111100011101",
                             6277 when "01111100011110",
                             6276 when "01111100011111",
                             6275 when "01111100100000",
                             6274 when "01111100100001",
                             6274 when "01111100100010",
                             6273 when "01111100100011",
                             6272 when "01111100100100",
                             6271 when "01111100100101",
                             6270 when "01111100100110",
                             6270 when "01111100100111",
                             6269 when "01111100101000",
                             6268 when "01111100101001",
                             6267 when "01111100101010",
                             6266 when "01111100101011",
                             6266 when "01111100101100",
                             6265 when "01111100101101",
                             6264 when "01111100101110",
                             6263 when "01111100101111",
                             6263 when "01111100110000",
                             6262 when "01111100110001",
                             6261 when "01111100110010",
                             6260 when "01111100110011",
                             6259 when "01111100110100",
                             6259 when "01111100110101",
                             6258 when "01111100110110",
                             6257 when "01111100110111",
                             6256 when "01111100111000",
                             6255 when "01111100111001",
                             6255 when "01111100111010",
                             6254 when "01111100111011",
                             6253 when "01111100111100",
                             6252 when "01111100111101",
                             6252 when "01111100111110",
                             6251 when "01111100111111",
                             6250 when "01111101000000",
                             6249 when "01111101000001",
                             6248 when "01111101000010",
                             6248 when "01111101000011",
                             6247 when "01111101000100",
                             6246 when "01111101000101",
                             6245 when "01111101000110",
                             6245 when "01111101000111",
                             6244 when "01111101001000",
                             6243 when "01111101001001",
                             6242 when "01111101001010",
                             6241 when "01111101001011",
                             6241 when "01111101001100",
                             6240 when "01111101001101",
                             6239 when "01111101001110",
                             6238 when "01111101001111",
                             6238 when "01111101010000",
                             6237 when "01111101010001",
                             6236 when "01111101010010",
                             6235 when "01111101010011",
                             6234 when "01111101010100",
                             6234 when "01111101010101",
                             6233 when "01111101010110",
                             6232 when "01111101010111",
                             6231 when "01111101011000",
                             6231 when "01111101011001",
                             6230 when "01111101011010",
                             6229 when "01111101011011",
                             6228 when "01111101011100",
                             6227 when "01111101011101",
                             6227 when "01111101011110",
                             6226 when "01111101011111",
                             6225 when "01111101100000",
                             6224 when "01111101100001",
                             6224 when "01111101100010",
                             6223 when "01111101100011",
                             6222 when "01111101100100",
                             6221 when "01111101100101",
                             6220 when "01111101100110",
                             6220 when "01111101100111",
                             6219 when "01111101101000",
                             6218 when "01111101101001",
                             6217 when "01111101101010",
                             6217 when "01111101101011",
                             6216 when "01111101101100",
                             6215 when "01111101101101",
                             6214 when "01111101101110",
                             6213 when "01111101101111",
                             6213 when "01111101110000",
                             6212 when "01111101110001",
                             6211 when "01111101110010",
                             6210 when "01111101110011",
                             6210 when "01111101110100",
                             6209 when "01111101110101",
                             6208 when "01111101110110",
                             6207 when "01111101110111",
                             6207 when "01111101111000",
                             6206 when "01111101111001",
                             6205 when "01111101111010",
                             6204 when "01111101111011",
                             6203 when "01111101111100",
                             6203 when "01111101111101",
                             6202 when "01111101111110",
                             6201 when "01111101111111",
                             6200 when "01111110000000",
                             6200 when "01111110000001",
                             6199 when "01111110000010",
                             6198 when "01111110000011",
                             6197 when "01111110000100",
                             6197 when "01111110000101",
                             6196 when "01111110000110",
                             6195 when "01111110000111",
                             6194 when "01111110001000",
                             6193 when "01111110001001",
                             6193 when "01111110001010",
                             6192 when "01111110001011",
                             6191 when "01111110001100",
                             6190 when "01111110001101",
                             6190 when "01111110001110",
                             6189 when "01111110001111",
                             6188 when "01111110010000",
                             6187 when "01111110010001",
                             6187 when "01111110010010",
                             6186 when "01111110010011",
                             6185 when "01111110010100",
                             6184 when "01111110010101",
                             6184 when "01111110010110",
                             6183 when "01111110010111",
                             6182 when "01111110011000",
                             6181 when "01111110011001",
                             6180 when "01111110011010",
                             6180 when "01111110011011",
                             6179 when "01111110011100",
                             6178 when "01111110011101",
                             6177 when "01111110011110",
                             6177 when "01111110011111",
                             6176 when "01111110100000",
                             6175 when "01111110100001",
                             6174 when "01111110100010",
                             6174 when "01111110100011",
                             6173 when "01111110100100",
                             6172 when "01111110100101",
                             6171 when "01111110100110",
                             6171 when "01111110100111",
                             6170 when "01111110101000",
                             6169 when "01111110101001",
                             6168 when "01111110101010",
                             6168 when "01111110101011",
                             6167 when "01111110101100",
                             6166 when "01111110101101",
                             6165 when "01111110101110",
                             6164 when "01111110101111",
                             6164 when "01111110110000",
                             6163 when "01111110110001",
                             6162 when "01111110110010",
                             6161 when "01111110110011",
                             6161 when "01111110110100",
                             6160 when "01111110110101",
                             6159 when "01111110110110",
                             6158 when "01111110110111",
                             6158 when "01111110111000",
                             6157 when "01111110111001",
                             6156 when "01111110111010",
                             6155 when "01111110111011",
                             6155 when "01111110111100",
                             6154 when "01111110111101",
                             6153 when "01111110111110",
                             6152 when "01111110111111",
                             6152 when "01111111000000",
                             6151 when "01111111000001",
                             6150 when "01111111000010",
                             6149 when "01111111000011",
                             6149 when "01111111000100",
                             6148 when "01111111000101",
                             6147 when "01111111000110",
                             6146 when "01111111000111",
                             6146 when "01111111001000",
                             6145 when "01111111001001",
                             6144 when "01111111001010",
                             6143 when "01111111001011",
                             6143 when "01111111001100",
                             6142 when "01111111001101",
                             6141 when "01111111001110",
                             6140 when "01111111001111",
                             6139 when "01111111010000",
                             6139 when "01111111010001",
                             6138 when "01111111010010",
                             6137 when "01111111010011",
                             6136 when "01111111010100",
                             6136 when "01111111010101",
                             6135 when "01111111010110",
                             6134 when "01111111010111",
                             6133 when "01111111011000",
                             6133 when "01111111011001",
                             6132 when "01111111011010",
                             6131 when "01111111011011",
                             6130 when "01111111011100",
                             6130 when "01111111011101",
                             6129 when "01111111011110",
                             6128 when "01111111011111",
                             6127 when "01111111100000",
                             6127 when "01111111100001",
                             6126 when "01111111100010",
                             6125 when "01111111100011",
                             6124 when "01111111100100",
                             6124 when "01111111100101",
                             6123 when "01111111100110",
                             6122 when "01111111100111",
                             6121 when "01111111101000",
                             6121 when "01111111101001",
                             6120 when "01111111101010",
                             6119 when "01111111101011",
                             6118 when "01111111101100",
                             6118 when "01111111101101",
                             6117 when "01111111101110",
                             6116 when "01111111101111",
                             6115 when "01111111110000",
                             6115 when "01111111110001",
                             6114 when "01111111110010",
                             6113 when "01111111110011",
                             6112 when "01111111110100",
                             6112 when "01111111110101",
                             6111 when "01111111110110",
                             6110 when "01111111110111",
                             6109 when "01111111111000",
                             6109 when "01111111111001",
                             6108 when "01111111111010",
                             6107 when "01111111111011",
                             6106 when "01111111111100",
                             6106 when "01111111111101",
                             6105 when "01111111111110",
                             6104 when "01111111111111",
                             6104 when "10000000000000",
                             6103 when "10000000000001",
                             6102 when "10000000000010",
                             6101 when "10000000000011",
                             6101 when "10000000000100",
                             6100 when "10000000000101",
                             6099 when "10000000000110",
                             6098 when "10000000000111",
                             6098 when "10000000001000",
                             6097 when "10000000001001",
                             6096 when "10000000001010",
                             6095 when "10000000001011",
                             6095 when "10000000001100",
                             6094 when "10000000001101",
                             6093 when "10000000001110",
                             6092 when "10000000001111",
                             6092 when "10000000010000",
                             6091 when "10000000010001",
                             6090 when "10000000010010",
                             6089 when "10000000010011",
                             6089 when "10000000010100",
                             6088 when "10000000010101",
                             6087 when "10000000010110",
                             6086 when "10000000010111",
                             6086 when "10000000011000",
                             6085 when "10000000011001",
                             6084 when "10000000011010",
                             6083 when "10000000011011",
                             6083 when "10000000011100",
                             6082 when "10000000011101",
                             6081 when "10000000011110",
                             6081 when "10000000011111",
                             6080 when "10000000100000",
                             6079 when "10000000100001",
                             6078 when "10000000100010",
                             6078 when "10000000100011",
                             6077 when "10000000100100",
                             6076 when "10000000100101",
                             6075 when "10000000100110",
                             6075 when "10000000100111",
                             6074 when "10000000101000",
                             6073 when "10000000101001",
                             6072 when "10000000101010",
                             6072 when "10000000101011",
                             6071 when "10000000101100",
                             6070 when "10000000101101",
                             6069 when "10000000101110",
                             6069 when "10000000101111",
                             6068 when "10000000110000",
                             6067 when "10000000110001",
                             6066 when "10000000110010",
                             6066 when "10000000110011",
                             6065 when "10000000110100",
                             6064 when "10000000110101",
                             6064 when "10000000110110",
                             6063 when "10000000110111",
                             6062 when "10000000111000",
                             6061 when "10000000111001",
                             6061 when "10000000111010",
                             6060 when "10000000111011",
                             6059 when "10000000111100",
                             6058 when "10000000111101",
                             6058 when "10000000111110",
                             6057 when "10000000111111",
                             6056 when "10000001000000",
                             6055 when "10000001000001",
                             6055 when "10000001000010",
                             6054 when "10000001000011",
                             6053 when "10000001000100",
                             6053 when "10000001000101",
                             6052 when "10000001000110",
                             6051 when "10000001000111",
                             6050 when "10000001001000",
                             6050 when "10000001001001",
                             6049 when "10000001001010",
                             6048 when "10000001001011",
                             6047 when "10000001001100",
                             6047 when "10000001001101",
                             6046 when "10000001001110",
                             6045 when "10000001001111",
                             6044 when "10000001010000",
                             6044 when "10000001010001",
                             6043 when "10000001010010",
                             6042 when "10000001010011",
                             6042 when "10000001010100",
                             6041 when "10000001010101",
                             6040 when "10000001010110",
                             6039 when "10000001010111",
                             6039 when "10000001011000",
                             6038 when "10000001011001",
                             6037 when "10000001011010",
                             6036 when "10000001011011",
                             6036 when "10000001011100",
                             6035 when "10000001011101",
                             6034 when "10000001011110",
                             6034 when "10000001011111",
                             6033 when "10000001100000",
                             6032 when "10000001100001",
                             6031 when "10000001100010",
                             6031 when "10000001100011",
                             6030 when "10000001100100",
                             6029 when "10000001100101",
                             6028 when "10000001100110",
                             6028 when "10000001100111",
                             6027 when "10000001101000",
                             6026 when "10000001101001",
                             6026 when "10000001101010",
                             6025 when "10000001101011",
                             6024 when "10000001101100",
                             6023 when "10000001101101",
                             6023 when "10000001101110",
                             6022 when "10000001101111",
                             6021 when "10000001110000",
                             6020 when "10000001110001",
                             6020 when "10000001110010",
                             6019 when "10000001110011",
                             6018 when "10000001110100",
                             6018 when "10000001110101",
                             6017 when "10000001110110",
                             6016 when "10000001110111",
                             6015 when "10000001111000",
                             6015 when "10000001111001",
                             6014 when "10000001111010",
                             6013 when "10000001111011",
                             6013 when "10000001111100",
                             6012 when "10000001111101",
                             6011 when "10000001111110",
                             6010 when "10000001111111",
                             6010 when "10000010000000",
                             6009 when "10000010000001",
                             6008 when "10000010000010",
                             6007 when "10000010000011",
                             6007 when "10000010000100",
                             6006 when "10000010000101",
                             6005 when "10000010000110",
                             6005 when "10000010000111",
                             6004 when "10000010001000",
                             6003 when "10000010001001",
                             6002 when "10000010001010",
                             6002 when "10000010001011",
                             6001 when "10000010001100",
                             6000 when "10000010001101",
                             6000 when "10000010001110",
                             5999 when "10000010001111",
                             5998 when "10000010010000",
                             5997 when "10000010010001",
                             5997 when "10000010010010",
                             5996 when "10000010010011",
                             5995 when "10000010010100",
                             5994 when "10000010010101",
                             5994 when "10000010010110",
                             5993 when "10000010010111",
                             5992 when "10000010011000",
                             5992 when "10000010011001",
                             5991 when "10000010011010",
                             5990 when "10000010011011",
                             5989 when "10000010011100",
                             5989 when "10000010011101",
                             5988 when "10000010011110",
                             5987 when "10000010011111",
                             5987 when "10000010100000",
                             5986 when "10000010100001",
                             5985 when "10000010100010",
                             5984 when "10000010100011",
                             5984 when "10000010100100",
                             5983 when "10000010100101",
                             5982 when "10000010100110",
                             5982 when "10000010100111",
                             5981 when "10000010101000",
                             5980 when "10000010101001",
                             5979 when "10000010101010",
                             5979 when "10000010101011",
                             5978 when "10000010101100",
                             5977 when "10000010101101",
                             5977 when "10000010101110",
                             5976 when "10000010101111",
                             5975 when "10000010110000",
                             5974 when "10000010110001",
                             5974 when "10000010110010",
                             5973 when "10000010110011",
                             5972 when "10000010110100",
                             5972 when "10000010110101",
                             5971 when "10000010110110",
                             5970 when "10000010110111",
                             5969 when "10000010111000",
                             5969 when "10000010111001",
                             5968 when "10000010111010",
                             5967 when "10000010111011",
                             5967 when "10000010111100",
                             5966 when "10000010111101",
                             5965 when "10000010111110",
                             5964 when "10000010111111",
                             5964 when "10000011000000",
                             5963 when "10000011000001",
                             5962 when "10000011000010",
                             5962 when "10000011000011",
                             5961 when "10000011000100",
                             5960 when "10000011000101",
                             5959 when "10000011000110",
                             5959 when "10000011000111",
                             5958 when "10000011001000",
                             5957 when "10000011001001",
                             5957 when "10000011001010",
                             5956 when "10000011001011",
                             5955 when "10000011001100",
                             5955 when "10000011001101",
                             5954 when "10000011001110",
                             5953 when "10000011001111",
                             5952 when "10000011010000",
                             5952 when "10000011010001",
                             5951 when "10000011010010",
                             5950 when "10000011010011",
                             5950 when "10000011010100",
                             5949 when "10000011010101",
                             5948 when "10000011010110",
                             5947 when "10000011010111",
                             5947 when "10000011011000",
                             5946 when "10000011011001",
                             5945 when "10000011011010",
                             5945 when "10000011011011",
                             5944 when "10000011011100",
                             5943 when "10000011011101",
                             5942 when "10000011011110",
                             5942 when "10000011011111",
                             5941 when "10000011100000",
                             5940 when "10000011100001",
                             5940 when "10000011100010",
                             5939 when "10000011100011",
                             5938 when "10000011100100",
                             5938 when "10000011100101",
                             5937 when "10000011100110",
                             5936 when "10000011100111",
                             5935 when "10000011101000",
                             5935 when "10000011101001",
                             5934 when "10000011101010",
                             5933 when "10000011101011",
                             5933 when "10000011101100",
                             5932 when "10000011101101",
                             5931 when "10000011101110",
                             5930 when "10000011101111",
                             5930 when "10000011110000",
                             5929 when "10000011110001",
                             5928 when "10000011110010",
                             5928 when "10000011110011",
                             5927 when "10000011110100",
                             5926 when "10000011110101",
                             5926 when "10000011110110",
                             5925 when "10000011110111",
                             5924 when "10000011111000",
                             5923 when "10000011111001",
                             5923 when "10000011111010",
                             5922 when "10000011111011",
                             5921 when "10000011111100",
                             5921 when "10000011111101",
                             5920 when "10000011111110",
                             5919 when "10000011111111",
                             5919 when "10000100000000",
                             5918 when "10000100000001",
                             5917 when "10000100000010",
                             5916 when "10000100000011",
                             5916 when "10000100000100",
                             5915 when "10000100000101",
                             5914 when "10000100000110",
                             5914 when "10000100000111",
                             5913 when "10000100001000",
                             5912 when "10000100001001",
                             5912 when "10000100001010",
                             5911 when "10000100001011",
                             5910 when "10000100001100",
                             5909 when "10000100001101",
                             5909 when "10000100001110",
                             5908 when "10000100001111",
                             5907 when "10000100010000",
                             5907 when "10000100010001",
                             5906 when "10000100010010",
                             5905 when "10000100010011",
                             5905 when "10000100010100",
                             5904 when "10000100010101",
                             5903 when "10000100010110",
                             5902 when "10000100010111",
                             5902 when "10000100011000",
                             5901 when "10000100011001",
                             5900 when "10000100011010",
                             5900 when "10000100011011",
                             5899 when "10000100011100",
                             5898 when "10000100011101",
                             5898 when "10000100011110",
                             5897 when "10000100011111",
                             5896 when "10000100100000",
                             5896 when "10000100100001",
                             5895 when "10000100100010",
                             5894 when "10000100100011",
                             5893 when "10000100100100",
                             5893 when "10000100100101",
                             5892 when "10000100100110",
                             5891 when "10000100100111",
                             5891 when "10000100101000",
                             5890 when "10000100101001",
                             5889 when "10000100101010",
                             5889 when "10000100101011",
                             5888 when "10000100101100",
                             5887 when "10000100101101",
                             5887 when "10000100101110",
                             5886 when "10000100101111",
                             5885 when "10000100110000",
                             5884 when "10000100110001",
                             5884 when "10000100110010",
                             5883 when "10000100110011",
                             5882 when "10000100110100",
                             5882 when "10000100110101",
                             5881 when "10000100110110",
                             5880 when "10000100110111",
                             5880 when "10000100111000",
                             5879 when "10000100111001",
                             5878 when "10000100111010",
                             5878 when "10000100111011",
                             5877 when "10000100111100",
                             5876 when "10000100111101",
                             5875 when "10000100111110",
                             5875 when "10000100111111",
                             5874 when "10000101000000",
                             5873 when "10000101000001",
                             5873 when "10000101000010",
                             5872 when "10000101000011",
                             5871 when "10000101000100",
                             5871 when "10000101000101",
                             5870 when "10000101000110",
                             5869 when "10000101000111",
                             5869 when "10000101001000",
                             5868 when "10000101001001",
                             5867 when "10000101001010",
                             5866 when "10000101001011",
                             5866 when "10000101001100",
                             5865 when "10000101001101",
                             5864 when "10000101001110",
                             5864 when "10000101001111",
                             5863 when "10000101010000",
                             5862 when "10000101010001",
                             5862 when "10000101010010",
                             5861 when "10000101010011",
                             5860 when "10000101010100",
                             5860 when "10000101010101",
                             5859 when "10000101010110",
                             5858 when "10000101010111",
                             5858 when "10000101011000",
                             5857 when "10000101011001",
                             5856 when "10000101011010",
                             5855 when "10000101011011",
                             5855 when "10000101011100",
                             5854 when "10000101011101",
                             5853 when "10000101011110",
                             5853 when "10000101011111",
                             5852 when "10000101100000",
                             5851 when "10000101100001",
                             5851 when "10000101100010",
                             5850 when "10000101100011",
                             5849 when "10000101100100",
                             5849 when "10000101100101",
                             5848 when "10000101100110",
                             5847 when "10000101100111",
                             5847 when "10000101101000",
                             5846 when "10000101101001",
                             5845 when "10000101101010",
                             5845 when "10000101101011",
                             5844 when "10000101101100",
                             5843 when "10000101101101",
                             5842 when "10000101101110",
                             5842 when "10000101101111",
                             5841 when "10000101110000",
                             5840 when "10000101110001",
                             5840 when "10000101110010",
                             5839 when "10000101110011",
                             5838 when "10000101110100",
                             5838 when "10000101110101",
                             5837 when "10000101110110",
                             5836 when "10000101110111",
                             5836 when "10000101111000",
                             5835 when "10000101111001",
                             5834 when "10000101111010",
                             5834 when "10000101111011",
                             5833 when "10000101111100",
                             5832 when "10000101111101",
                             5832 when "10000101111110",
                             5831 when "10000101111111",
                             5830 when "10000110000000",
                             5830 when "10000110000001",
                             5829 when "10000110000010",
                             5828 when "10000110000011",
                             5828 when "10000110000100",
                             5827 when "10000110000101",
                             5826 when "10000110000110",
                             5825 when "10000110000111",
                             5825 when "10000110001000",
                             5824 when "10000110001001",
                             5823 when "10000110001010",
                             5823 when "10000110001011",
                             5822 when "10000110001100",
                             5821 when "10000110001101",
                             5821 when "10000110001110",
                             5820 when "10000110001111",
                             5819 when "10000110010000",
                             5819 when "10000110010001",
                             5818 when "10000110010010",
                             5817 when "10000110010011",
                             5817 when "10000110010100",
                             5816 when "10000110010101",
                             5815 when "10000110010110",
                             5815 when "10000110010111",
                             5814 when "10000110011000",
                             5813 when "10000110011001",
                             5813 when "10000110011010",
                             5812 when "10000110011011",
                             5811 when "10000110011100",
                             5811 when "10000110011101",
                             5810 when "10000110011110",
                             5809 when "10000110011111",
                             5809 when "10000110100000",
                             5808 when "10000110100001",
                             5807 when "10000110100010",
                             5807 when "10000110100011",
                             5806 when "10000110100100",
                             5805 when "10000110100101",
                             5805 when "10000110100110",
                             5804 when "10000110100111",
                             5803 when "10000110101000",
                             5802 when "10000110101001",
                             5802 when "10000110101010",
                             5801 when "10000110101011",
                             5800 when "10000110101100",
                             5800 when "10000110101101",
                             5799 when "10000110101110",
                             5798 when "10000110101111",
                             5798 when "10000110110000",
                             5797 when "10000110110001",
                             5796 when "10000110110010",
                             5796 when "10000110110011",
                             5795 when "10000110110100",
                             5794 when "10000110110101",
                             5794 when "10000110110110",
                             5793 when "10000110110111",
                             5792 when "10000110111000",
                             5792 when "10000110111001",
                             5791 when "10000110111010",
                             5790 when "10000110111011",
                             5790 when "10000110111100",
                             5789 when "10000110111101",
                             5788 when "10000110111110",
                             5788 when "10000110111111",
                             5787 when "10000111000000",
                             5786 when "10000111000001",
                             5786 when "10000111000010",
                             5785 when "10000111000011",
                             5784 when "10000111000100",
                             5784 when "10000111000101",
                             5783 when "10000111000110",
                             5782 when "10000111000111",
                             5782 when "10000111001000",
                             5781 when "10000111001001",
                             5780 when "10000111001010",
                             5780 when "10000111001011",
                             5779 when "10000111001100",
                             5778 when "10000111001101",
                             5778 when "10000111001110",
                             5777 when "10000111001111",
                             5776 when "10000111010000",
                             5776 when "10000111010001",
                             5775 when "10000111010010",
                             5774 when "10000111010011",
                             5774 when "10000111010100",
                             5773 when "10000111010101",
                             5772 when "10000111010110",
                             5772 when "10000111010111",
                             5771 when "10000111011000",
                             5770 when "10000111011001",
                             5770 when "10000111011010",
                             5769 when "10000111011011",
                             5768 when "10000111011100",
                             5768 when "10000111011101",
                             5767 when "10000111011110",
                             5766 when "10000111011111",
                             5766 when "10000111100000",
                             5765 when "10000111100001",
                             5764 when "10000111100010",
                             5764 when "10000111100011",
                             5763 when "10000111100100",
                             5762 when "10000111100101",
                             5762 when "10000111100110",
                             5761 when "10000111100111",
                             5760 when "10000111101000",
                             5760 when "10000111101001",
                             5759 when "10000111101010",
                             5758 when "10000111101011",
                             5758 when "10000111101100",
                             5757 when "10000111101101",
                             5756 when "10000111101110",
                             5756 when "10000111101111",
                             5755 when "10000111110000",
                             5754 when "10000111110001",
                             5754 when "10000111110010",
                             5753 when "10000111110011",
                             5752 when "10000111110100",
                             5752 when "10000111110101",
                             5751 when "10000111110110",
                             5750 when "10000111110111",
                             5750 when "10000111111000",
                             5749 when "10000111111001",
                             5748 when "10000111111010",
                             5748 when "10000111111011",
                             5747 when "10000111111100",
                             5746 when "10000111111101",
                             5746 when "10000111111110",
                             5745 when "10000111111111",
                             5744 when "10001000000000",
                             5744 when "10001000000001",
                             5743 when "10001000000010",
                             5743 when "10001000000011",
                             5742 when "10001000000100",
                             5741 when "10001000000101",
                             5741 when "10001000000110",
                             5740 when "10001000000111",
                             5739 when "10001000001000",
                             5739 when "10001000001001",
                             5738 when "10001000001010",
                             5737 when "10001000001011",
                             5737 when "10001000001100",
                             5736 when "10001000001101",
                             5735 when "10001000001110",
                             5735 when "10001000001111",
                             5734 when "10001000010000",
                             5733 when "10001000010001",
                             5733 when "10001000010010",
                             5732 when "10001000010011",
                             5731 when "10001000010100",
                             5731 when "10001000010101",
                             5730 when "10001000010110",
                             5729 when "10001000010111",
                             5729 when "10001000011000",
                             5728 when "10001000011001",
                             5727 when "10001000011010",
                             5727 when "10001000011011",
                             5726 when "10001000011100",
                             5725 when "10001000011101",
                             5725 when "10001000011110",
                             5724 when "10001000011111",
                             5723 when "10001000100000",
                             5723 when "10001000100001",
                             5722 when "10001000100010",
                             5721 when "10001000100011",
                             5721 when "10001000100100",
                             5720 when "10001000100101",
                             5720 when "10001000100110",
                             5719 when "10001000100111",
                             5718 when "10001000101000",
                             5718 when "10001000101001",
                             5717 when "10001000101010",
                             5716 when "10001000101011",
                             5716 when "10001000101100",
                             5715 when "10001000101101",
                             5714 when "10001000101110",
                             5714 when "10001000101111",
                             5713 when "10001000110000",
                             5712 when "10001000110001",
                             5712 when "10001000110010",
                             5711 when "10001000110011",
                             5710 when "10001000110100",
                             5710 when "10001000110101",
                             5709 when "10001000110110",
                             5708 when "10001000110111",
                             5708 when "10001000111000",
                             5707 when "10001000111001",
                             5706 when "10001000111010",
                             5706 when "10001000111011",
                             5705 when "10001000111100",
                             5705 when "10001000111101",
                             5704 when "10001000111110",
                             5703 when "10001000111111",
                             5703 when "10001001000000",
                             5702 when "10001001000001",
                             5701 when "10001001000010",
                             5701 when "10001001000011",
                             5700 when "10001001000100",
                             5699 when "10001001000101",
                             5699 when "10001001000110",
                             5698 when "10001001000111",
                             5697 when "10001001001000",
                             5697 when "10001001001001",
                             5696 when "10001001001010",
                             5695 when "10001001001011",
                             5695 when "10001001001100",
                             5694 when "10001001001101",
                             5693 when "10001001001110",
                             5693 when "10001001001111",
                             5692 when "10001001010000",
                             5692 when "10001001010001",
                             5691 when "10001001010010",
                             5690 when "10001001010011",
                             5690 when "10001001010100",
                             5689 when "10001001010101",
                             5688 when "10001001010110",
                             5688 when "10001001010111",
                             5687 when "10001001011000",
                             5686 when "10001001011001",
                             5686 when "10001001011010",
                             5685 when "10001001011011",
                             5684 when "10001001011100",
                             5684 when "10001001011101",
                             5683 when "10001001011110",
                             5682 when "10001001011111",
                             5682 when "10001001100000",
                             5681 when "10001001100001",
                             5681 when "10001001100010",
                             5680 when "10001001100011",
                             5679 when "10001001100100",
                             5679 when "10001001100101",
                             5678 when "10001001100110",
                             5677 when "10001001100111",
                             5677 when "10001001101000",
                             5676 when "10001001101001",
                             5675 when "10001001101010",
                             5675 when "10001001101011",
                             5674 when "10001001101100",
                             5673 when "10001001101101",
                             5673 when "10001001101110",
                             5672 when "10001001101111",
                             5672 when "10001001110000",
                             5671 when "10001001110001",
                             5670 when "10001001110010",
                             5670 when "10001001110011",
                             5669 when "10001001110100",
                             5668 when "10001001110101",
                             5668 when "10001001110110",
                             5667 when "10001001110111",
                             5666 when "10001001111000",
                             5666 when "10001001111001",
                             5665 when "10001001111010",
                             5664 when "10001001111011",
                             5664 when "10001001111100",
                             5663 when "10001001111101",
                             5663 when "10001001111110",
                             5662 when "10001001111111",
                             5661 when "10001010000000",
                             5661 when "10001010000001",
                             5660 when "10001010000010",
                             5659 when "10001010000011",
                             5659 when "10001010000100",
                             5658 when "10001010000101",
                             5657 when "10001010000110",
                             5657 when "10001010000111",
                             5656 when "10001010001000",
                             5655 when "10001010001001",
                             5655 when "10001010001010",
                             5654 when "10001010001011",
                             5654 when "10001010001100",
                             5653 when "10001010001101",
                             5652 when "10001010001110",
                             5652 when "10001010001111",
                             5651 when "10001010010000",
                             5650 when "10001010010001",
                             5650 when "10001010010010",
                             5649 when "10001010010011",
                             5648 when "10001010010100",
                             5648 when "10001010010101",
                             5647 when "10001010010110",
                             5647 when "10001010010111",
                             5646 when "10001010011000",
                             5645 when "10001010011001",
                             5645 when "10001010011010",
                             5644 when "10001010011011",
                             5643 when "10001010011100",
                             5643 when "10001010011101",
                             5642 when "10001010011110",
                             5641 when "10001010011111",
                             5641 when "10001010100000",
                             5640 when "10001010100001",
                             5640 when "10001010100010",
                             5639 when "10001010100011",
                             5638 when "10001010100100",
                             5638 when "10001010100101",
                             5637 when "10001010100110",
                             5636 when "10001010100111",
                             5636 when "10001010101000",
                             5635 when "10001010101001",
                             5634 when "10001010101010",
                             5634 when "10001010101011",
                             5633 when "10001010101100",
                             5633 when "10001010101101",
                             5632 when "10001010101110",
                             5631 when "10001010101111",
                             5631 when "10001010110000",
                             5630 when "10001010110001",
                             5629 when "10001010110010",
                             5629 when "10001010110011",
                             5628 when "10001010110100",
                             5627 when "10001010110101",
                             5627 when "10001010110110",
                             5626 when "10001010110111",
                             5626 when "10001010111000",
                             5625 when "10001010111001",
                             5624 when "10001010111010",
                             5624 when "10001010111011",
                             5623 when "10001010111100",
                             5622 when "10001010111101",
                             5622 when "10001010111110",
                             5621 when "10001010111111",
                             5621 when "10001011000000",
                             5620 when "10001011000001",
                             5619 when "10001011000010",
                             5619 when "10001011000011",
                             5618 when "10001011000100",
                             5617 when "10001011000101",
                             5617 when "10001011000110",
                             5616 when "10001011000111",
                             5615 when "10001011001000",
                             5615 when "10001011001001",
                             5614 when "10001011001010",
                             5614 when "10001011001011",
                             5613 when "10001011001100",
                             5612 when "10001011001101",
                             5612 when "10001011001110",
                             5611 when "10001011001111",
                             5610 when "10001011010000",
                             5610 when "10001011010001",
                             5609 when "10001011010010",
                             5609 when "10001011010011",
                             5608 when "10001011010100",
                             5607 when "10001011010101",
                             5607 when "10001011010110",
                             5606 when "10001011010111",
                             5605 when "10001011011000",
                             5605 when "10001011011001",
                             5604 when "10001011011010",
                             5603 when "10001011011011",
                             5603 when "10001011011100",
                             5602 when "10001011011101",
                             5602 when "10001011011110",
                             5601 when "10001011011111",
                             5600 when "10001011100000",
                             5600 when "10001011100001",
                             5599 when "10001011100010",
                             5598 when "10001011100011",
                             5598 when "10001011100100",
                             5597 when "10001011100101",
                             5597 when "10001011100110",
                             5596 when "10001011100111",
                             5595 when "10001011101000",
                             5595 when "10001011101001",
                             5594 when "10001011101010",
                             5593 when "10001011101011",
                             5593 when "10001011101100",
                             5592 when "10001011101101",
                             5592 when "10001011101110",
                             5591 when "10001011101111",
                             5590 when "10001011110000",
                             5590 when "10001011110001",
                             5589 when "10001011110010",
                             5588 when "10001011110011",
                             5588 when "10001011110100",
                             5587 when "10001011110101",
                             5587 when "10001011110110",
                             5586 when "10001011110111",
                             5585 when "10001011111000",
                             5585 when "10001011111001",
                             5584 when "10001011111010",
                             5583 when "10001011111011",
                             5583 when "10001011111100",
                             5582 when "10001011111101",
                             5582 when "10001011111110",
                             5581 when "10001011111111",
                             5580 when "10001100000000",
                             5580 when "10001100000001",
                             5579 when "10001100000010",
                             5578 when "10001100000011",
                             5578 when "10001100000100",
                             5577 when "10001100000101",
                             5577 when "10001100000110",
                             5576 when "10001100000111",
                             5575 when "10001100001000",
                             5575 when "10001100001001",
                             5574 when "10001100001010",
                             5574 when "10001100001011",
                             5573 when "10001100001100",
                             5572 when "10001100001101",
                             5572 when "10001100001110",
                             5571 when "10001100001111",
                             5570 when "10001100010000",
                             5570 when "10001100010001",
                             5569 when "10001100010010",
                             5569 when "10001100010011",
                             5568 when "10001100010100",
                             5567 when "10001100010101",
                             5567 when "10001100010110",
                             5566 when "10001100010111",
                             5565 when "10001100011000",
                             5565 when "10001100011001",
                             5564 when "10001100011010",
                             5564 when "10001100011011",
                             5563 when "10001100011100",
                             5562 when "10001100011101",
                             5562 when "10001100011110",
                             5561 when "10001100011111",
                             5560 when "10001100100000",
                             5560 when "10001100100001",
                             5559 when "10001100100010",
                             5559 when "10001100100011",
                             5558 when "10001100100100",
                             5557 when "10001100100101",
                             5557 when "10001100100110",
                             5556 when "10001100100111",
                             5556 when "10001100101000",
                             5555 when "10001100101001",
                             5554 when "10001100101010",
                             5554 when "10001100101011",
                             5553 when "10001100101100",
                             5552 when "10001100101101",
                             5552 when "10001100101110",
                             5551 when "10001100101111",
                             5551 when "10001100110000",
                             5550 when "10001100110001",
                             5549 when "10001100110010",
                             5549 when "10001100110011",
                             5548 when "10001100110100",
                             5548 when "10001100110101",
                             5547 when "10001100110110",
                             5546 when "10001100110111",
                             5546 when "10001100111000",
                             5545 when "10001100111001",
                             5544 when "10001100111010",
                             5544 when "10001100111011",
                             5543 when "10001100111100",
                             5543 when "10001100111101",
                             5542 when "10001100111110",
                             5541 when "10001100111111",
                             5541 when "10001101000000",
                             5540 when "10001101000001",
                             5540 when "10001101000010",
                             5539 when "10001101000011",
                             5538 when "10001101000100",
                             5538 when "10001101000101",
                             5537 when "10001101000110",
                             5536 when "10001101000111",
                             5536 when "10001101001000",
                             5535 when "10001101001001",
                             5535 when "10001101001010",
                             5534 when "10001101001011",
                             5533 when "10001101001100",
                             5533 when "10001101001101",
                             5532 when "10001101001110",
                             5532 when "10001101001111",
                             5531 when "10001101010000",
                             5530 when "10001101010001",
                             5530 when "10001101010010",
                             5529 when "10001101010011",
                             5529 when "10001101010100",
                             5528 when "10001101010101",
                             5527 when "10001101010110",
                             5527 when "10001101010111",
                             5526 when "10001101011000",
                             5525 when "10001101011001",
                             5525 when "10001101011010",
                             5524 when "10001101011011",
                             5524 when "10001101011100",
                             5523 when "10001101011101",
                             5522 when "10001101011110",
                             5522 when "10001101011111",
                             5521 when "10001101100000",
                             5521 when "10001101100001",
                             5520 when "10001101100010",
                             5519 when "10001101100011",
                             5519 when "10001101100100",
                             5518 when "10001101100101",
                             5518 when "10001101100110",
                             5517 when "10001101100111",
                             5516 when "10001101101000",
                             5516 when "10001101101001",
                             5515 when "10001101101010",
                             5515 when "10001101101011",
                             5514 when "10001101101100",
                             5513 when "10001101101101",
                             5513 when "10001101101110",
                             5512 when "10001101101111",
                             5511 when "10001101110000",
                             5511 when "10001101110001",
                             5510 when "10001101110010",
                             5510 when "10001101110011",
                             5509 when "10001101110100",
                             5508 when "10001101110101",
                             5508 when "10001101110110",
                             5507 when "10001101110111",
                             5507 when "10001101111000",
                             5506 when "10001101111001",
                             5505 when "10001101111010",
                             5505 when "10001101111011",
                             5504 when "10001101111100",
                             5504 when "10001101111101",
                             5503 when "10001101111110",
                             5502 when "10001101111111",
                             5502 when "10001110000000",
                             5501 when "10001110000001",
                             5501 when "10001110000010",
                             5500 when "10001110000011",
                             5499 when "10001110000100",
                             5499 when "10001110000101",
                             5498 when "10001110000110",
                             5498 when "10001110000111",
                             5497 when "10001110001000",
                             5496 when "10001110001001",
                             5496 when "10001110001010",
                             5495 when "10001110001011",
                             5495 when "10001110001100",
                             5494 when "10001110001101",
                             5493 when "10001110001110",
                             5493 when "10001110001111",
                             5492 when "10001110010000",
                             5491 when "10001110010001",
                             5491 when "10001110010010",
                             5490 when "10001110010011",
                             5490 when "10001110010100",
                             5489 when "10001110010101",
                             5488 when "10001110010110",
                             5488 when "10001110010111",
                             5487 when "10001110011000",
                             5487 when "10001110011001",
                             5486 when "10001110011010",
                             5485 when "10001110011011",
                             5485 when "10001110011100",
                             5484 when "10001110011101",
                             5484 when "10001110011110",
                             5483 when "10001110011111",
                             5482 when "10001110100000",
                             5482 when "10001110100001",
                             5481 when "10001110100010",
                             5481 when "10001110100011",
                             5480 when "10001110100100",
                             5479 when "10001110100101",
                             5479 when "10001110100110",
                             5478 when "10001110100111",
                             5478 when "10001110101000",
                             5477 when "10001110101001",
                             5476 when "10001110101010",
                             5476 when "10001110101011",
                             5475 when "10001110101100",
                             5475 when "10001110101101",
                             5474 when "10001110101110",
                             5473 when "10001110101111",
                             5473 when "10001110110000",
                             5472 when "10001110110001",
                             5472 when "10001110110010",
                             5471 when "10001110110011",
                             5470 when "10001110110100",
                             5470 when "10001110110101",
                             5469 when "10001110110110",
                             5469 when "10001110110111",
                             5468 when "10001110111000",
                             5467 when "10001110111001",
                             5467 when "10001110111010",
                             5466 when "10001110111011",
                             5466 when "10001110111100",
                             5465 when "10001110111101",
                             5464 when "10001110111110",
                             5464 when "10001110111111",
                             5463 when "10001111000000",
                             5463 when "10001111000001",
                             5462 when "10001111000010",
                             5461 when "10001111000011",
                             5461 when "10001111000100",
                             5460 when "10001111000101",
                             5460 when "10001111000110",
                             5459 when "10001111000111",
                             5459 when "10001111001000",
                             5458 when "10001111001001",
                             5457 when "10001111001010",
                             5457 when "10001111001011",
                             5456 when "10001111001100",
                             5456 when "10001111001101",
                             5455 when "10001111001110",
                             5454 when "10001111001111",
                             5454 when "10001111010000",
                             5453 when "10001111010001",
                             5453 when "10001111010010",
                             5452 when "10001111010011",
                             5451 when "10001111010100",
                             5451 when "10001111010101",
                             5450 when "10001111010110",
                             5450 when "10001111010111",
                             5449 when "10001111011000",
                             5448 when "10001111011001",
                             5448 when "10001111011010",
                             5447 when "10001111011011",
                             5447 when "10001111011100",
                             5446 when "10001111011101",
                             5445 when "10001111011110",
                             5445 when "10001111011111",
                             5444 when "10001111100000",
                             5444 when "10001111100001",
                             5443 when "10001111100010",
                             5442 when "10001111100011",
                             5442 when "10001111100100",
                             5441 when "10001111100101",
                             5441 when "10001111100110",
                             5440 when "10001111100111",
                             5440 when "10001111101000",
                             5439 when "10001111101001",
                             5438 when "10001111101010",
                             5438 when "10001111101011",
                             5437 when "10001111101100",
                             5437 when "10001111101101",
                             5436 when "10001111101110",
                             5435 when "10001111101111",
                             5435 when "10001111110000",
                             5434 when "10001111110001",
                             5434 when "10001111110010",
                             5433 when "10001111110011",
                             5432 when "10001111110100",
                             5432 when "10001111110101",
                             5431 when "10001111110110",
                             5431 when "10001111110111",
                             5430 when "10001111111000",
                             5429 when "10001111111001",
                             5429 when "10001111111010",
                             5428 when "10001111111011",
                             5428 when "10001111111100",
                             5427 when "10001111111101",
                             5427 when "10001111111110",
                             5426 when "10001111111111",
                             5425 when "10010000000000",
                             5425 when "10010000000001",
                             5424 when "10010000000010",
                             5424 when "10010000000011",
                             5423 when "10010000000100",
                             5422 when "10010000000101",
                             5422 when "10010000000110",
                             5421 when "10010000000111",
                             5421 when "10010000001000",
                             5420 when "10010000001001",
                             5419 when "10010000001010",
                             5419 when "10010000001011",
                             5418 when "10010000001100",
                             5418 when "10010000001101",
                             5417 when "10010000001110",
                             5417 when "10010000001111",
                             5416 when "10010000010000",
                             5415 when "10010000010001",
                             5415 when "10010000010010",
                             5414 when "10010000010011",
                             5414 when "10010000010100",
                             5413 when "10010000010101",
                             5412 when "10010000010110",
                             5412 when "10010000010111",
                             5411 when "10010000011000",
                             5411 when "10010000011001",
                             5410 when "10010000011010",
                             5409 when "10010000011011",
                             5409 when "10010000011100",
                             5408 when "10010000011101",
                             5408 when "10010000011110",
                             5407 when "10010000011111",
                             5407 when "10010000100000",
                             5406 when "10010000100001",
                             5405 when "10010000100010",
                             5405 when "10010000100011",
                             5404 when "10010000100100",
                             5404 when "10010000100101",
                             5403 when "10010000100110",
                             5402 when "10010000100111",
                             5402 when "10010000101000",
                             5401 when "10010000101001",
                             5401 when "10010000101010",
                             5400 when "10010000101011",
                             5400 when "10010000101100",
                             5399 when "10010000101101",
                             5398 when "10010000101110",
                             5398 when "10010000101111",
                             5397 when "10010000110000",
                             5397 when "10010000110001",
                             5396 when "10010000110010",
                             5395 when "10010000110011",
                             5395 when "10010000110100",
                             5394 when "10010000110101",
                             5394 when "10010000110110",
                             5393 when "10010000110111",
                             5393 when "10010000111000",
                             5392 when "10010000111001",
                             5391 when "10010000111010",
                             5391 when "10010000111011",
                             5390 when "10010000111100",
                             5390 when "10010000111101",
                             5389 when "10010000111110",
                             5389 when "10010000111111",
                             5388 when "10010001000000",
                             5387 when "10010001000001",
                             5387 when "10010001000010",
                             5386 when "10010001000011",
                             5386 when "10010001000100",
                             5385 when "10010001000101",
                             5384 when "10010001000110",
                             5384 when "10010001000111",
                             5383 when "10010001001000",
                             5383 when "10010001001001",
                             5382 when "10010001001010",
                             5382 when "10010001001011",
                             5381 when "10010001001100",
                             5380 when "10010001001101",
                             5380 when "10010001001110",
                             5379 when "10010001001111",
                             5379 when "10010001010000",
                             5378 when "10010001010001",
                             5378 when "10010001010010",
                             5377 when "10010001010011",
                             5376 when "10010001010100",
                             5376 when "10010001010101",
                             5375 when "10010001010110",
                             5375 when "10010001010111",
                             5374 when "10010001011000",
                             5373 when "10010001011001",
                             5373 when "10010001011010",
                             5372 when "10010001011011",
                             5372 when "10010001011100",
                             5371 when "10010001011101",
                             5371 when "10010001011110",
                             5370 when "10010001011111",
                             5369 when "10010001100000",
                             5369 when "10010001100001",
                             5368 when "10010001100010",
                             5368 when "10010001100011",
                             5367 when "10010001100100",
                             5367 when "10010001100101",
                             5366 when "10010001100110",
                             5365 when "10010001100111",
                             5365 when "10010001101000",
                             5364 when "10010001101001",
                             5364 when "10010001101010",
                             5363 when "10010001101011",
                             5363 when "10010001101100",
                             5362 when "10010001101101",
                             5361 when "10010001101110",
                             5361 when "10010001101111",
                             5360 when "10010001110000",
                             5360 when "10010001110001",
                             5359 when "10010001110010",
                             5358 when "10010001110011",
                             5358 when "10010001110100",
                             5357 when "10010001110101",
                             5357 when "10010001110110",
                             5356 when "10010001110111",
                             5356 when "10010001111000",
                             5355 when "10010001111001",
                             5354 when "10010001111010",
                             5354 when "10010001111011",
                             5353 when "10010001111100",
                             5353 when "10010001111101",
                             5352 when "10010001111110",
                             5352 when "10010001111111",
                             5351 when "10010010000000",
                             5350 when "10010010000001",
                             5350 when "10010010000010",
                             5349 when "10010010000011",
                             5349 when "10010010000100",
                             5348 when "10010010000101",
                             5348 when "10010010000110",
                             5347 when "10010010000111",
                             5346 when "10010010001000",
                             5346 when "10010010001001",
                             5345 when "10010010001010",
                             5345 when "10010010001011",
                             5344 when "10010010001100",
                             5344 when "10010010001101",
                             5343 when "10010010001110",
                             5342 when "10010010001111",
                             5342 when "10010010010000",
                             5341 when "10010010010001",
                             5341 when "10010010010010",
                             5340 when "10010010010011",
                             5340 when "10010010010100",
                             5339 when "10010010010101",
                             5338 when "10010010010110",
                             5338 when "10010010010111",
                             5337 when "10010010011000",
                             5337 when "10010010011001",
                             5336 when "10010010011010",
                             5336 when "10010010011011",
                             5335 when "10010010011100",
                             5334 when "10010010011101",
                             5334 when "10010010011110",
                             5333 when "10010010011111",
                             5333 when "10010010100000",
                             5332 when "10010010100001",
                             5332 when "10010010100010",
                             5331 when "10010010100011",
                             5330 when "10010010100100",
                             5330 when "10010010100101",
                             5329 when "10010010100110",
                             5329 when "10010010100111",
                             5328 when "10010010101000",
                             5328 when "10010010101001",
                             5327 when "10010010101010",
                             5327 when "10010010101011",
                             5326 when "10010010101100",
                             5325 when "10010010101101",
                             5325 when "10010010101110",
                             5324 when "10010010101111",
                             5324 when "10010010110000",
                             5323 when "10010010110001",
                             5323 when "10010010110010",
                             5322 when "10010010110011",
                             5321 when "10010010110100",
                             5321 when "10010010110101",
                             5320 when "10010010110110",
                             5320 when "10010010110111",
                             5319 when "10010010111000",
                             5319 when "10010010111001",
                             5318 when "10010010111010",
                             5317 when "10010010111011",
                             5317 when "10010010111100",
                             5316 when "10010010111101",
                             5316 when "10010010111110",
                             5315 when "10010010111111",
                             5315 when "10010011000000",
                             5314 when "10010011000001",
                             5313 when "10010011000010",
                             5313 when "10010011000011",
                             5312 when "10010011000100",
                             5312 when "10010011000101",
                             5311 when "10010011000110",
                             5311 when "10010011000111",
                             5310 when "10010011001000",
                             5310 when "10010011001001",
                             5309 when "10010011001010",
                             5308 when "10010011001011",
                             5308 when "10010011001100",
                             5307 when "10010011001101",
                             5307 when "10010011001110",
                             5306 when "10010011001111",
                             5306 when "10010011010000",
                             5305 when "10010011010001",
                             5304 when "10010011010010",
                             5304 when "10010011010011",
                             5303 when "10010011010100",
                             5303 when "10010011010101",
                             5302 when "10010011010110",
                             5302 when "10010011010111",
                             5301 when "10010011011000",
                             5301 when "10010011011001",
                             5300 when "10010011011010",
                             5299 when "10010011011011",
                             5299 when "10010011011100",
                             5298 when "10010011011101",
                             5298 when "10010011011110",
                             5297 when "10010011011111",
                             5297 when "10010011100000",
                             5296 when "10010011100001",
                             5295 when "10010011100010",
                             5295 when "10010011100011",
                             5294 when "10010011100100",
                             5294 when "10010011100101",
                             5293 when "10010011100110",
                             5293 when "10010011100111",
                             5292 when "10010011101000",
                             5292 when "10010011101001",
                             5291 when "10010011101010",
                             5290 when "10010011101011",
                             5290 when "10010011101100",
                             5289 when "10010011101101",
                             5289 when "10010011101110",
                             5288 when "10010011101111",
                             5288 when "10010011110000",
                             5287 when "10010011110001",
                             5287 when "10010011110010",
                             5286 when "10010011110011",
                             5285 when "10010011110100",
                             5285 when "10010011110101",
                             5284 when "10010011110110",
                             5284 when "10010011110111",
                             5283 when "10010011111000",
                             5283 when "10010011111001",
                             5282 when "10010011111010",
                             5282 when "10010011111011",
                             5281 when "10010011111100",
                             5280 when "10010011111101",
                             5280 when "10010011111110",
                             5279 when "10010011111111",
                             5279 when "10010100000000",
                             5278 when "10010100000001",
                             5278 when "10010100000010",
                             5277 when "10010100000011",
                             5276 when "10010100000100",
                             5276 when "10010100000101",
                             5275 when "10010100000110",
                             5275 when "10010100000111",
                             5274 when "10010100001000",
                             5274 when "10010100001001",
                             5273 when "10010100001010",
                             5273 when "10010100001011",
                             5272 when "10010100001100",
                             5271 when "10010100001101",
                             5271 when "10010100001110",
                             5270 when "10010100001111",
                             5270 when "10010100010000",
                             5269 when "10010100010001",
                             5269 when "10010100010010",
                             5268 when "10010100010011",
                             5268 when "10010100010100",
                             5267 when "10010100010101",
                             5266 when "10010100010110",
                             5266 when "10010100010111",
                             5265 when "10010100011000",
                             5265 when "10010100011001",
                             5264 when "10010100011010",
                             5264 when "10010100011011",
                             5263 when "10010100011100",
                             5263 when "10010100011101",
                             5262 when "10010100011110",
                             5261 when "10010100011111",
                             5261 when "10010100100000",
                             5260 when "10010100100001",
                             5260 when "10010100100010",
                             5259 when "10010100100011",
                             5259 when "10010100100100",
                             5258 when "10010100100101",
                             5258 when "10010100100110",
                             5257 when "10010100100111",
                             5257 when "10010100101000",
                             5256 when "10010100101001",
                             5255 when "10010100101010",
                             5255 when "10010100101011",
                             5254 when "10010100101100",
                             5254 when "10010100101101",
                             5253 when "10010100101110",
                             5253 when "10010100101111",
                             5252 when "10010100110000",
                             5252 when "10010100110001",
                             5251 when "10010100110010",
                             5250 when "10010100110011",
                             5250 when "10010100110100",
                             5249 when "10010100110101",
                             5249 when "10010100110110",
                             5248 when "10010100110111",
                             5248 when "10010100111000",
                             5247 when "10010100111001",
                             5247 when "10010100111010",
                             5246 when "10010100111011",
                             5245 when "10010100111100",
                             5245 when "10010100111101",
                             5244 when "10010100111110",
                             5244 when "10010100111111",
                             5243 when "10010101000000",
                             5243 when "10010101000001",
                             5242 when "10010101000010",
                             5242 when "10010101000011",
                             5241 when "10010101000100",
                             5241 when "10010101000101",
                             5240 when "10010101000110",
                             5239 when "10010101000111",
                             5239 when "10010101001000",
                             5238 when "10010101001001",
                             5238 when "10010101001010",
                             5237 when "10010101001011",
                             5237 when "10010101001100",
                             5236 when "10010101001101",
                             5236 when "10010101001110",
                             5235 when "10010101001111",
                             5235 when "10010101010000",
                             5234 when "10010101010001",
                             5233 when "10010101010010",
                             5233 when "10010101010011",
                             5232 when "10010101010100",
                             5232 when "10010101010101",
                             5231 when "10010101010110",
                             5231 when "10010101010111",
                             5230 when "10010101011000",
                             5230 when "10010101011001",
                             5229 when "10010101011010",
                             5228 when "10010101011011",
                             5228 when "10010101011100",
                             5227 when "10010101011101",
                             5227 when "10010101011110",
                             5226 when "10010101011111",
                             5226 when "10010101100000",
                             5225 when "10010101100001",
                             5225 when "10010101100010",
                             5224 when "10010101100011",
                             5224 when "10010101100100",
                             5223 when "10010101100101",
                             5222 when "10010101100110",
                             5222 when "10010101100111",
                             5221 when "10010101101000",
                             5221 when "10010101101001",
                             5220 when "10010101101010",
                             5220 when "10010101101011",
                             5219 when "10010101101100",
                             5219 when "10010101101101",
                             5218 when "10010101101110",
                             5218 when "10010101101111",
                             5217 when "10010101110000",
                             5216 when "10010101110001",
                             5216 when "10010101110010",
                             5215 when "10010101110011",
                             5215 when "10010101110100",
                             5214 when "10010101110101",
                             5214 when "10010101110110",
                             5213 when "10010101110111",
                             5213 when "10010101111000",
                             5212 when "10010101111001",
                             5212 when "10010101111010",
                             5211 when "10010101111011",
                             5211 when "10010101111100",
                             5210 when "10010101111101",
                             5209 when "10010101111110",
                             5209 when "10010101111111",
                             5208 when "10010110000000",
                             5208 when "10010110000001",
                             5207 when "10010110000010",
                             5207 when "10010110000011",
                             5206 when "10010110000100",
                             5206 when "10010110000101",
                             5205 when "10010110000110",
                             5205 when "10010110000111",
                             5204 when "10010110001000",
                             5203 when "10010110001001",
                             5203 when "10010110001010",
                             5202 when "10010110001011",
                             5202 when "10010110001100",
                             5201 when "10010110001101",
                             5201 when "10010110001110",
                             5200 when "10010110001111",
                             5200 when "10010110010000",
                             5199 when "10010110010001",
                             5199 when "10010110010010",
                             5198 when "10010110010011",
                             5198 when "10010110010100",
                             5197 when "10010110010101",
                             5196 when "10010110010110",
                             5196 when "10010110010111",
                             5195 when "10010110011000",
                             5195 when "10010110011001",
                             5194 when "10010110011010",
                             5194 when "10010110011011",
                             5193 when "10010110011100",
                             5193 when "10010110011101",
                             5192 when "10010110011110",
                             5192 when "10010110011111",
                             5191 when "10010110100000",
                             5190 when "10010110100001",
                             5190 when "10010110100010",
                             5189 when "10010110100011",
                             5189 when "10010110100100",
                             5188 when "10010110100101",
                             5188 when "10010110100110",
                             5187 when "10010110100111",
                             5187 when "10010110101000",
                             5186 when "10010110101001",
                             5186 when "10010110101010",
                             5185 when "10010110101011",
                             5185 when "10010110101100",
                             5184 when "10010110101101",
                             5183 when "10010110101110",
                             5183 when "10010110101111",
                             5182 when "10010110110000",
                             5182 when "10010110110001",
                             5181 when "10010110110010",
                             5181 when "10010110110011",
                             5180 when "10010110110100",
                             5180 when "10010110110101",
                             5179 when "10010110110110",
                             5179 when "10010110110111",
                             5178 when "10010110111000",
                             5178 when "10010110111001",
                             5177 when "10010110111010",
                             5177 when "10010110111011",
                             5176 when "10010110111100",
                             5175 when "10010110111101",
                             5175 when "10010110111110",
                             5174 when "10010110111111",
                             5174 when "10010111000000",
                             5173 when "10010111000001",
                             5173 when "10010111000010",
                             5172 when "10010111000011",
                             5172 when "10010111000100",
                             5171 when "10010111000101",
                             5171 when "10010111000110",
                             5170 when "10010111000111",
                             5170 when "10010111001000",
                             5169 when "10010111001001",
                             5168 when "10010111001010",
                             5168 when "10010111001011",
                             5167 when "10010111001100",
                             5167 when "10010111001101",
                             5166 when "10010111001110",
                             5166 when "10010111001111",
                             5165 when "10010111010000",
                             5165 when "10010111010001",
                             5164 when "10010111010010",
                             5164 when "10010111010011",
                             5163 when "10010111010100",
                             5163 when "10010111010101",
                             5162 when "10010111010110",
                             5162 when "10010111010111",
                             5161 when "10010111011000",
                             5160 when "10010111011001",
                             5160 when "10010111011010",
                             5159 when "10010111011011",
                             5159 when "10010111011100",
                             5158 when "10010111011101",
                             5158 when "10010111011110",
                             5157 when "10010111011111",
                             5157 when "10010111100000",
                             5156 when "10010111100001",
                             5156 when "10010111100010",
                             5155 when "10010111100011",
                             5155 when "10010111100100",
                             5154 when "10010111100101",
                             5154 when "10010111100110",
                             5153 when "10010111100111",
                             5153 when "10010111101000",
                             5152 when "10010111101001",
                             5151 when "10010111101010",
                             5151 when "10010111101011",
                             5150 when "10010111101100",
                             5150 when "10010111101101",
                             5149 when "10010111101110",
                             5149 when "10010111101111",
                             5148 when "10010111110000",
                             5148 when "10010111110001",
                             5147 when "10010111110010",
                             5147 when "10010111110011",
                             5146 when "10010111110100",
                             5146 when "10010111110101",
                             5145 when "10010111110110",
                             5145 when "10010111110111",
                             5144 when "10010111111000",
                             5144 when "10010111111001",
                             5143 when "10010111111010",
                             5142 when "10010111111011",
                             5142 when "10010111111100",
                             5141 when "10010111111101",
                             5141 when "10010111111110",
                             5140 when "10010111111111",
                             5140 when "10011000000000",
                             5139 when "10011000000001",
                             5139 when "10011000000010",
                             5138 when "10011000000011",
                             5138 when "10011000000100",
                             5137 when "10011000000101",
                             5137 when "10011000000110",
                             5136 when "10011000000111",
                             5136 when "10011000001000",
                             5135 when "10011000001001",
                             5135 when "10011000001010",
                             5134 when "10011000001011",
                             5133 when "10011000001100",
                             5133 when "10011000001101",
                             5132 when "10011000001110",
                             5132 when "10011000001111",
                             5131 when "10011000010000",
                             5131 when "10011000010001",
                             5130 when "10011000010010",
                             5130 when "10011000010011",
                             5129 when "10011000010100",
                             5129 when "10011000010101",
                             5128 when "10011000010110",
                             5128 when "10011000010111",
                             5127 when "10011000011000",
                             5127 when "10011000011001",
                             5126 when "10011000011010",
                             5126 when "10011000011011",
                             5125 when "10011000011100",
                             5125 when "10011000011101",
                             5124 when "10011000011110",
                             5123 when "10011000011111",
                             5123 when "10011000100000",
                             5122 when "10011000100001",
                             5122 when "10011000100010",
                             5121 when "10011000100011",
                             5121 when "10011000100100",
                             5120 when "10011000100101",
                             5120 when "10011000100110",
                             5119 when "10011000100111",
                             5119 when "10011000101000",
                             5118 when "10011000101001",
                             5118 when "10011000101010",
                             5117 when "10011000101011",
                             5117 when "10011000101100",
                             5116 when "10011000101101",
                             5116 when "10011000101110",
                             5115 when "10011000101111",
                             5115 when "10011000110000",
                             5114 when "10011000110001",
                             5114 when "10011000110010",
                             5113 when "10011000110011",
                             5112 when "10011000110100",
                             5112 when "10011000110101",
                             5111 when "10011000110110",
                             5111 when "10011000110111",
                             5110 when "10011000111000",
                             5110 when "10011000111001",
                             5109 when "10011000111010",
                             5109 when "10011000111011",
                             5108 when "10011000111100",
                             5108 when "10011000111101",
                             5107 when "10011000111110",
                             5107 when "10011000111111",
                             5106 when "10011001000000",
                             5106 when "10011001000001",
                             5105 when "10011001000010",
                             5105 when "10011001000011",
                             5104 when "10011001000100",
                             5104 when "10011001000101",
                             5103 when "10011001000110",
                             5103 when "10011001000111",
                             5102 when "10011001001000",
                             5102 when "10011001001001",
                             5101 when "10011001001010",
                             5100 when "10011001001011",
                             5100 when "10011001001100",
                             5099 when "10011001001101",
                             5099 when "10011001001110",
                             5098 when "10011001001111",
                             5098 when "10011001010000",
                             5097 when "10011001010001",
                             5097 when "10011001010010",
                             5096 when "10011001010011",
                             5096 when "10011001010100",
                             5095 when "10011001010101",
                             5095 when "10011001010110",
                             5094 when "10011001010111",
                             5094 when "10011001011000",
                             5093 when "10011001011001",
                             5093 when "10011001011010",
                             5092 when "10011001011011",
                             5092 when "10011001011100",
                             5091 when "10011001011101",
                             5091 when "10011001011110",
                             5090 when "10011001011111",
                             5090 when "10011001100000",
                             5089 when "10011001100001",
                             5089 when "10011001100010",
                             5088 when "10011001100011",
                             5088 when "10011001100100",
                             5087 when "10011001100101",
                             5086 when "10011001100110",
                             5086 when "10011001100111",
                             5085 when "10011001101000",
                             5085 when "10011001101001",
                             5084 when "10011001101010",
                             5084 when "10011001101011",
                             5083 when "10011001101100",
                             5083 when "10011001101101",
                             5082 when "10011001101110",
                             5082 when "10011001101111",
                             5081 when "10011001110000",
                             5081 when "10011001110001",
                             5080 when "10011001110010",
                             5080 when "10011001110011",
                             5079 when "10011001110100",
                             5079 when "10011001110101",
                             5078 when "10011001110110",
                             5078 when "10011001110111",
                             5077 when "10011001111000",
                             5077 when "10011001111001",
                             5076 when "10011001111010",
                             5076 when "10011001111011",
                             5075 when "10011001111100",
                             5075 when "10011001111101",
                             5074 when "10011001111110",
                             5074 when "10011001111111",
                             5073 when "10011010000000",
                             5073 when "10011010000001",
                             5072 when "10011010000010",
                             5072 when "10011010000011",
                             5071 when "10011010000100",
                             5070 when "10011010000101",
                             5070 when "10011010000110",
                             5069 when "10011010000111",
                             5069 when "10011010001000",
                             5068 when "10011010001001",
                             5068 when "10011010001010",
                             5067 when "10011010001011",
                             5067 when "10011010001100",
                             5066 when "10011010001101",
                             5066 when "10011010001110",
                             5065 when "10011010001111",
                             5065 when "10011010010000",
                             5064 when "10011010010001",
                             5064 when "10011010010010",
                             5063 when "10011010010011",
                             5063 when "10011010010100",
                             5062 when "10011010010101",
                             5062 when "10011010010110",
                             5061 when "10011010010111",
                             5061 when "10011010011000",
                             5060 when "10011010011001",
                             5060 when "10011010011010",
                             5059 when "10011010011011",
                             5059 when "10011010011100",
                             5058 when "10011010011101",
                             5058 when "10011010011110",
                             5057 when "10011010011111",
                             5057 when "10011010100000",
                             5056 when "10011010100001",
                             5056 when "10011010100010",
                             5055 when "10011010100011",
                             5055 when "10011010100100",
                             5054 when "10011010100101",
                             5054 when "10011010100110",
                             5053 when "10011010100111",
                             5053 when "10011010101000",
                             5052 when "10011010101001",
                             5052 when "10011010101010",
                             5051 when "10011010101011",
                             5051 when "10011010101100",
                             5050 when "10011010101101",
                             5049 when "10011010101110",
                             5049 when "10011010101111",
                             5048 when "10011010110000",
                             5048 when "10011010110001",
                             5047 when "10011010110010",
                             5047 when "10011010110011",
                             5046 when "10011010110100",
                             5046 when "10011010110101",
                             5045 when "10011010110110",
                             5045 when "10011010110111",
                             5044 when "10011010111000",
                             5044 when "10011010111001",
                             5043 when "10011010111010",
                             5043 when "10011010111011",
                             5042 when "10011010111100",
                             5042 when "10011010111101",
                             5041 when "10011010111110",
                             5041 when "10011010111111",
                             5040 when "10011011000000",
                             5040 when "10011011000001",
                             5039 when "10011011000010",
                             5039 when "10011011000011",
                             5038 when "10011011000100",
                             5038 when "10011011000101",
                             5037 when "10011011000110",
                             5037 when "10011011000111",
                             5036 when "10011011001000",
                             5036 when "10011011001001",
                             5035 when "10011011001010",
                             5035 when "10011011001011",
                             5034 when "10011011001100",
                             5034 when "10011011001101",
                             5033 when "10011011001110",
                             5033 when "10011011001111",
                             5032 when "10011011010000",
                             5032 when "10011011010001",
                             5031 when "10011011010010",
                             5031 when "10011011010011",
                             5030 when "10011011010100",
                             5030 when "10011011010101",
                             5029 when "10011011010110",
                             5029 when "10011011010111",
                             5028 when "10011011011000",
                             5028 when "10011011011001",
                             5027 when "10011011011010",
                             5027 when "10011011011011",
                             5026 when "10011011011100",
                             5026 when "10011011011101",
                             5025 when "10011011011110",
                             5025 when "10011011011111",
                             5024 when "10011011100000",
                             5024 when "10011011100001",
                             5023 when "10011011100010",
                             5023 when "10011011100011",
                             5022 when "10011011100100",
                             5022 when "10011011100101",
                             5021 when "10011011100110",
                             5021 when "10011011100111",
                             5020 when "10011011101000",
                             5020 when "10011011101001",
                             5019 when "10011011101010",
                             5019 when "10011011101011",
                             5018 when "10011011101100",
                             5018 when "10011011101101",
                             5017 when "10011011101110",
                             5017 when "10011011101111",
                             5016 when "10011011110000",
                             5016 when "10011011110001",
                             5015 when "10011011110010",
                             5015 when "10011011110011",
                             5014 when "10011011110100",
                             5014 when "10011011110101",
                             5013 when "10011011110110",
                             5013 when "10011011110111",
                             5012 when "10011011111000",
                             5012 when "10011011111001",
                             5011 when "10011011111010",
                             5011 when "10011011111011",
                             5010 when "10011011111100",
                             5010 when "10011011111101",
                             5009 when "10011011111110",
                             5009 when "10011011111111",
                             5008 when "10011100000000",
                             5008 when "10011100000001",
                             5007 when "10011100000010",
                             5007 when "10011100000011",
                             5006 when "10011100000100",
                             5006 when "10011100000101",
                             5005 when "10011100000110",
                             5005 when "10011100000111",
                             5004 when "10011100001000",
                             5004 when "10011100001001",
                             5003 when "10011100001010",
                             5003 when "10011100001011",
                             5002 when "10011100001100",
                             5002 when "10011100001101",
                             5001 when "10011100001110",
                             5001 when "10011100001111",
                             5000 when "10011100010000",
                             5000 when "10011100010001",
                             4999 when "10011100010010",
                             4999 when "10011100010011",
                             4998 when "10011100010100",
                             4998 when "10011100010101",
                             4997 when "10011100010110",
                             4997 when "10011100010111",
                             4996 when "10011100011000",
                             4996 when "10011100011001",
                             4995 when "10011100011010",
                             4995 when "10011100011011",
                             4994 when "10011100011100",
                             4994 when "10011100011101",
                             4993 when "10011100011110",
                             4993 when "10011100011111",
                             4992 when "10011100100000",
                             4992 when "10011100100001",
                             4991 when "10011100100010",
                             4991 when "10011100100011",
                             4990 when "10011100100100",
                             4990 when "10011100100101",
                             4989 when "10011100100110",
                             4989 when "10011100100111",
                             4988 when "10011100101000",
                             4988 when "10011100101001",
                             4987 when "10011100101010",
                             4987 when "10011100101011",
                             4986 when "10011100101100",
                             4986 when "10011100101101",
                             4985 when "10011100101110",
                             4985 when "10011100101111",
                             4984 when "10011100110000",
                             4984 when "10011100110001",
                             4983 when "10011100110010",
                             4983 when "10011100110011",
                             4982 when "10011100110100",
                             4982 when "10011100110101",
                             4981 when "10011100110110",
                             4981 when "10011100110111",
                             4980 when "10011100111000",
                             4980 when "10011100111001",
                             4979 when "10011100111010",
                             4979 when "10011100111011",
                             4978 when "10011100111100",
                             4978 when "10011100111101",
                             4977 when "10011100111110",
                             4977 when "10011100111111",
                             4976 when "10011101000000",
                             4976 when "10011101000001",
                             4975 when "10011101000010",
                             4975 when "10011101000011",
                             4974 when "10011101000100",
                             4974 when "10011101000101",
                             4973 when "10011101000110",
                             4973 when "10011101000111",
                             4972 when "10011101001000",
                             4972 when "10011101001001",
                             4971 when "10011101001010",
                             4971 when "10011101001011",
                             4970 when "10011101001100",
                             4970 when "10011101001101",
                             4969 when "10011101001110",
                             4969 when "10011101001111",
                             4968 when "10011101010000",
                             4968 when "10011101010001",
                             4967 when "10011101010010",
                             4967 when "10011101010011",
                             4966 when "10011101010100",
                             4966 when "10011101010101",
                             4965 when "10011101010110",
                             4965 when "10011101010111",
                             4964 when "10011101011000",
                             4964 when "10011101011001",
                             4963 when "10011101011010",
                             4963 when "10011101011011",
                             4962 when "10011101011100",
                             4962 when "10011101011101",
                             4961 when "10011101011110",
                             4961 when "10011101011111",
                             4960 when "10011101100000",
                             4960 when "10011101100001",
                             4959 when "10011101100010",
                             4959 when "10011101100011",
                             4958 when "10011101100100",
                             4958 when "10011101100101",
                             4957 when "10011101100110",
                             4957 when "10011101100111",
                             4956 when "10011101101000",
                             4956 when "10011101101001",
                             4955 when "10011101101010",
                             4955 when "10011101101011",
                             4954 when "10011101101100",
                             4954 when "10011101101101",
                             4953 when "10011101101110",
                             4953 when "10011101101111",
                             4952 when "10011101110000",
                             4952 when "10011101110001",
                             4951 when "10011101110010",
                             4951 when "10011101110011",
                             4950 when "10011101110100",
                             4950 when "10011101110101",
                             4950 when "10011101110110",
                             4949 when "10011101110111",
                             4949 when "10011101111000",
                             4948 when "10011101111001",
                             4948 when "10011101111010",
                             4947 when "10011101111011",
                             4947 when "10011101111100",
                             4946 when "10011101111101",
                             4946 when "10011101111110",
                             4945 when "10011101111111",
                             4945 when "10011110000000",
                             4944 when "10011110000001",
                             4944 when "10011110000010",
                             4943 when "10011110000011",
                             4943 when "10011110000100",
                             4942 when "10011110000101",
                             4942 when "10011110000110",
                             4941 when "10011110000111",
                             4941 when "10011110001000",
                             4940 when "10011110001001",
                             4940 when "10011110001010",
                             4939 when "10011110001011",
                             4939 when "10011110001100",
                             4938 when "10011110001101",
                             4938 when "10011110001110",
                             4937 when "10011110001111",
                             4937 when "10011110010000",
                             4936 when "10011110010001",
                             4936 when "10011110010010",
                             4935 when "10011110010011",
                             4935 when "10011110010100",
                             4934 when "10011110010101",
                             4934 when "10011110010110",
                             4933 when "10011110010111",
                             4933 when "10011110011000",
                             4932 when "10011110011001",
                             4932 when "10011110011010",
                             4931 when "10011110011011",
                             4931 when "10011110011100",
                             4930 when "10011110011101",
                             4930 when "10011110011110",
                             4930 when "10011110011111",
                             4929 when "10011110100000",
                             4929 when "10011110100001",
                             4928 when "10011110100010",
                             4928 when "10011110100011",
                             4927 when "10011110100100",
                             4927 when "10011110100101",
                             4926 when "10011110100110",
                             4926 when "10011110100111",
                             4925 when "10011110101000",
                             4925 when "10011110101001",
                             4924 when "10011110101010",
                             4924 when "10011110101011",
                             4923 when "10011110101100",
                             4923 when "10011110101101",
                             4922 when "10011110101110",
                             4922 when "10011110101111",
                             4921 when "10011110110000",
                             4921 when "10011110110001",
                             4920 when "10011110110010",
                             4920 when "10011110110011",
                             4919 when "10011110110100",
                             4919 when "10011110110101",
                             4918 when "10011110110110",
                             4918 when "10011110110111",
                             4917 when "10011110111000",
                             4917 when "10011110111001",
                             4916 when "10011110111010",
                             4916 when "10011110111011",
                             4915 when "10011110111100",
                             4915 when "10011110111101",
                             4914 when "10011110111110",
                             4914 when "10011110111111",
                             4914 when "10011111000000",
                             4913 when "10011111000001",
                             4913 when "10011111000010",
                             4912 when "10011111000011",
                             4912 when "10011111000100",
                             4911 when "10011111000101",
                             4911 when "10011111000110",
                             4910 when "10011111000111",
                             4910 when "10011111001000",
                             4909 when "10011111001001",
                             4909 when "10011111001010",
                             4908 when "10011111001011",
                             4908 when "10011111001100",
                             4907 when "10011111001101",
                             4907 when "10011111001110",
                             4906 when "10011111001111",
                             4906 when "10011111010000",
                             4905 when "10011111010001",
                             4905 when "10011111010010",
                             4904 when "10011111010011",
                             4904 when "10011111010100",
                             4903 when "10011111010101",
                             4903 when "10011111010110",
                             4902 when "10011111010111",
                             4902 when "10011111011000",
                             4901 when "10011111011001",
                             4901 when "10011111011010",
                             4901 when "10011111011011",
                             4900 when "10011111011100",
                             4900 when "10011111011101",
                             4899 when "10011111011110",
                             4899 when "10011111011111",
                             4898 when "10011111100000",
                             4898 when "10011111100001",
                             4897 when "10011111100010",
                             4897 when "10011111100011",
                             4896 when "10011111100100",
                             4896 when "10011111100101",
                             4895 when "10011111100110",
                             4895 when "10011111100111",
                             4894 when "10011111101000",
                             4894 when "10011111101001",
                             4893 when "10011111101010",
                             4893 when "10011111101011",
                             4892 when "10011111101100",
                             4892 when "10011111101101",
                             4891 when "10011111101110",
                             4891 when "10011111101111",
                             4890 when "10011111110000",
                             4890 when "10011111110001",
                             4889 when "10011111110010",
                             4889 when "10011111110011",
                             4889 when "10011111110100",
                             4888 when "10011111110101",
                             4888 when "10011111110110",
                             4887 when "10011111110111",
                             4887 when "10011111111000",
                             4886 when "10011111111001",
                             4886 when "10011111111010",
                             4885 when "10011111111011",
                             4885 when "10011111111100",
                             4884 when "10011111111101",
                             4884 when "10011111111110",
                             4883 when "10011111111111",
                             4883 when "10100000000000",
                             4882 when "10100000000001",
                             4882 when "10100000000010",
                             4881 when "10100000000011",
                             4881 when "10100000000100",
                             4880 when "10100000000101",
                             4880 when "10100000000110",
                             4879 when "10100000000111",
                             4879 when "10100000001000",
                             4879 when "10100000001001",
                             4878 when "10100000001010",
                             4878 when "10100000001011",
                             4877 when "10100000001100",
                             4877 when "10100000001101",
                             4876 when "10100000001110",
                             4876 when "10100000001111",
                             4875 when "10100000010000",
                             4875 when "10100000010001",
                             4874 when "10100000010010",
                             4874 when "10100000010011",
                             4873 when "10100000010100",
                             4873 when "10100000010101",
                             4872 when "10100000010110",
                             4872 when "10100000010111",
                             4871 when "10100000011000",
                             4871 when "10100000011001",
                             4870 when "10100000011010",
                             4870 when "10100000011011",
                             4869 when "10100000011100",
                             4869 when "10100000011101",
                             4869 when "10100000011110",
                             4868 when "10100000011111",
                             4868 when "10100000100000",
                             4867 when "10100000100001",
                             4867 when "10100000100010",
                             4866 when "10100000100011",
                             4866 when "10100000100100",
                             4865 when "10100000100101",
                             4865 when "10100000100110",
                             4864 when "10100000100111",
                             4864 when "10100000101000",
                             4863 when "10100000101001",
                             4863 when "10100000101010",
                             4862 when "10100000101011",
                             4862 when "10100000101100",
                             4861 when "10100000101101",
                             4861 when "10100000101110",
                             4861 when "10100000101111",
                             4860 when "10100000110000",
                             4860 when "10100000110001",
                             4859 when "10100000110010",
                             4859 when "10100000110011",
                             4858 when "10100000110100",
                             4858 when "10100000110101",
                             4857 when "10100000110110",
                             4857 when "10100000110111",
                             4856 when "10100000111000",
                             4856 when "10100000111001",
                             4855 when "10100000111010",
                             4855 when "10100000111011",
                             4854 when "10100000111100",
                             4854 when "10100000111101",
                             4853 when "10100000111110",
                             4853 when "10100000111111",
                             4852 when "10100001000000",
                             4852 when "10100001000001",
                             4852 when "10100001000010",
                             4851 when "10100001000011",
                             4851 when "10100001000100",
                             4850 when "10100001000101",
                             4850 when "10100001000110",
                             4849 when "10100001000111",
                             4849 when "10100001001000",
                             4848 when "10100001001001",
                             4848 when "10100001001010",
                             4847 when "10100001001011",
                             4847 when "10100001001100",
                             4846 when "10100001001101",
                             4846 when "10100001001110",
                             4845 when "10100001001111",
                             4845 when "10100001010000",
                             4844 when "10100001010001",
                             4844 when "10100001010010",
                             4844 when "10100001010011",
                             4843 when "10100001010100",
                             4843 when "10100001010101",
                             4842 when "10100001010110",
                             4842 when "10100001010111",
                             4841 when "10100001011000",
                             4841 when "10100001011001",
                             4840 when "10100001011010",
                             4840 when "10100001011011",
                             4839 when "10100001011100",
                             4839 when "10100001011101",
                             4838 when "10100001011110",
                             4838 when "10100001011111",
                             4837 when "10100001100000",
                             4837 when "10100001100001",
                             4837 when "10100001100010",
                             4836 when "10100001100011",
                             4836 when "10100001100100",
                             4835 when "10100001100101",
                             4835 when "10100001100110",
                             4834 when "10100001100111",
                             4834 when "10100001101000",
                             4833 when "10100001101001",
                             4833 when "10100001101010",
                             4832 when "10100001101011",
                             4832 when "10100001101100",
                             4831 when "10100001101101",
                             4831 when "10100001101110",
                             4830 when "10100001101111",
                             4830 when "10100001110000",
                             4830 when "10100001110001",
                             4829 when "10100001110010",
                             4829 when "10100001110011",
                             4828 when "10100001110100",
                             4828 when "10100001110101",
                             4827 when "10100001110110",
                             4827 when "10100001110111",
                             4826 when "10100001111000",
                             4826 when "10100001111001",
                             4825 when "10100001111010",
                             4825 when "10100001111011",
                             4824 when "10100001111100",
                             4824 when "10100001111101",
                             4823 when "10100001111110",
                             4823 when "10100001111111",
                             4823 when "10100010000000",
                             4822 when "10100010000001",
                             4822 when "10100010000010",
                             4821 when "10100010000011",
                             4821 when "10100010000100",
                             4820 when "10100010000101",
                             4820 when "10100010000110",
                             4819 when "10100010000111",
                             4819 when "10100010001000",
                             4818 when "10100010001001",
                             4818 when "10100010001010",
                             4817 when "10100010001011",
                             4817 when "10100010001100",
                             4816 when "10100010001101",
                             4816 when "10100010001110",
                             4816 when "10100010001111",
                             4815 when "10100010010000",
                             4815 when "10100010010001",
                             4814 when "10100010010010",
                             4814 when "10100010010011",
                             4813 when "10100010010100",
                             4813 when "10100010010101",
                             4812 when "10100010010110",
                             4812 when "10100010010111",
                             4811 when "10100010011000",
                             4811 when "10100010011001",
                             4810 when "10100010011010",
                             4810 when "10100010011011",
                             4810 when "10100010011100",
                             4809 when "10100010011101",
                             4809 when "10100010011110",
                             4808 when "10100010011111",
                             4808 when "10100010100000",
                             4807 when "10100010100001",
                             4807 when "10100010100010",
                             4806 when "10100010100011",
                             4806 when "10100010100100",
                             4805 when "10100010100101",
                             4805 when "10100010100110",
                             4804 when "10100010100111",
                             4804 when "10100010101000",
                             4804 when "10100010101001",
                             4803 when "10100010101010",
                             4803 when "10100010101011",
                             4802 when "10100010101100",
                             4802 when "10100010101101",
                             4801 when "10100010101110",
                             4801 when "10100010101111",
                             4800 when "10100010110000",
                             4800 when "10100010110001",
                             4799 when "10100010110010",
                             4799 when "10100010110011",
                             4798 when "10100010110100",
                             4798 when "10100010110101",
                             4798 when "10100010110110",
                             4797 when "10100010110111",
                             4797 when "10100010111000",
                             4796 when "10100010111001",
                             4796 when "10100010111010",
                             4795 when "10100010111011",
                             4795 when "10100010111100",
                             4794 when "10100010111101",
                             4794 when "10100010111110",
                             4793 when "10100010111111",
                             4793 when "10100011000000",
                             4792 when "10100011000001",
                             4792 when "10100011000010",
                             4792 when "10100011000011",
                             4791 when "10100011000100",
                             4791 when "10100011000101",
                             4790 when "10100011000110",
                             4790 when "10100011000111",
                             4789 when "10100011001000",
                             4789 when "10100011001001",
                             4788 when "10100011001010",
                             4788 when "10100011001011",
                             4787 when "10100011001100",
                             4787 when "10100011001101",
                             4787 when "10100011001110",
                             4786 when "10100011001111",
                             4786 when "10100011010000",
                             4785 when "10100011010001",
                             4785 when "10100011010010",
                             4784 when "10100011010011",
                             4784 when "10100011010100",
                             4783 when "10100011010101",
                             4783 when "10100011010110",
                             4782 when "10100011010111",
                             4782 when "10100011011000",
                             4781 when "10100011011001",
                             4781 when "10100011011010",
                             4781 when "10100011011011",
                             4780 when "10100011011100",
                             4780 when "10100011011101",
                             4779 when "10100011011110",
                             4779 when "10100011011111",
                             4778 when "10100011100000",
                             4778 when "10100011100001",
                             4777 when "10100011100010",
                             4777 when "10100011100011",
                             4776 when "10100011100100",
                             4776 when "10100011100101",
                             4776 when "10100011100110",
                             4775 when "10100011100111",
                             4775 when "10100011101000",
                             4774 when "10100011101001",
                             4774 when "10100011101010",
                             4773 when "10100011101011",
                             4773 when "10100011101100",
                             4772 when "10100011101101",
                             4772 when "10100011101110",
                             4771 when "10100011101111",
                             4771 when "10100011110000",
                             4771 when "10100011110001",
                             4770 when "10100011110010",
                             4770 when "10100011110011",
                             4769 when "10100011110100",
                             4769 when "10100011110101",
                             4768 when "10100011110110",
                             4768 when "10100011110111",
                             4767 when "10100011111000",
                             4767 when "10100011111001",
                             4766 when "10100011111010",
                             4766 when "10100011111011",
                             4766 when "10100011111100",
                             4765 when "10100011111101",
                             4765 when "10100011111110",
                             4764 when "10100011111111",
                             4764 when "10100100000000",
                             4763 when "10100100000001",
                             4763 when "10100100000010",
                             4762 when "10100100000011",
                             4762 when "10100100000100",
                             4761 when "10100100000101",
                             4761 when "10100100000110",
                             4761 when "10100100000111",
                             4760 when "10100100001000",
                             4760 when "10100100001001",
                             4759 when "10100100001010",
                             4759 when "10100100001011",
                             4758 when "10100100001100",
                             4758 when "10100100001101",
                             4757 when "10100100001110",
                             4757 when "10100100001111",
                             4756 when "10100100010000",
                             4756 when "10100100010001",
                             4756 when "10100100010010",
                             4755 when "10100100010011",
                             4755 when "10100100010100",
                             4754 when "10100100010101",
                             4754 when "10100100010110",
                             4753 when "10100100010111",
                             4753 when "10100100011000",
                             4752 when "10100100011001",
                             4752 when "10100100011010",
                             4751 when "10100100011011",
                             4751 when "10100100011100",
                             4751 when "10100100011101",
                             4750 when "10100100011110",
                             4750 when "10100100011111",
                             4749 when "10100100100000",
                             4749 when "10100100100001",
                             4748 when "10100100100010",
                             4748 when "10100100100011",
                             4747 when "10100100100100",
                             4747 when "10100100100101",
                             4747 when "10100100100110",
                             4746 when "10100100100111",
                             4746 when "10100100101000",
                             4745 when "10100100101001",
                             4745 when "10100100101010",
                             4744 when "10100100101011",
                             4744 when "10100100101100",
                             4743 when "10100100101101",
                             4743 when "10100100101110",
                             4742 when "10100100101111",
                             4742 when "10100100110000",
                             4742 when "10100100110001",
                             4741 when "10100100110010",
                             4741 when "10100100110011",
                             4740 when "10100100110100",
                             4740 when "10100100110101",
                             4739 when "10100100110110",
                             4739 when "10100100110111",
                             4738 when "10100100111000",
                             4738 when "10100100111001",
                             4738 when "10100100111010",
                             4737 when "10100100111011",
                             4737 when "10100100111100",
                             4736 when "10100100111101",
                             4736 when "10100100111110",
                             4735 when "10100100111111",
                             4735 when "10100101000000",
                             4734 when "10100101000001",
                             4734 when "10100101000010",
                             4734 when "10100101000011",
                             4733 when "10100101000100",
                             4733 when "10100101000101",
                             4732 when "10100101000110",
                             4732 when "10100101000111",
                             4731 when "10100101001000",
                             4731 when "10100101001001",
                             4730 when "10100101001010",
                             4730 when "10100101001011",
                             4729 when "10100101001100",
                             4729 when "10100101001101",
                             4729 when "10100101001110",
                             4728 when "10100101001111",
                             4728 when "10100101010000",
                             4727 when "10100101010001",
                             4727 when "10100101010010",
                             4726 when "10100101010011",
                             4726 when "10100101010100",
                             4725 when "10100101010101",
                             4725 when "10100101010110",
                             4725 when "10100101010111",
                             4724 when "10100101011000",
                             4724 when "10100101011001",
                             4723 when "10100101011010",
                             4723 when "10100101011011",
                             4722 when "10100101011100",
                             4722 when "10100101011101",
                             4721 when "10100101011110",
                             4721 when "10100101011111",
                             4721 when "10100101100000",
                             4720 when "10100101100001",
                             4720 when "10100101100010",
                             4719 when "10100101100011",
                             4719 when "10100101100100",
                             4718 when "10100101100101",
                             4718 when "10100101100110",
                             4717 when "10100101100111",
                             4717 when "10100101101000",
                             4717 when "10100101101001",
                             4716 when "10100101101010",
                             4716 when "10100101101011",
                             4715 when "10100101101100",
                             4715 when "10100101101101",
                             4714 when "10100101101110",
                             4714 when "10100101101111",
                             4713 when "10100101110000",
                             4713 when "10100101110001",
                             4713 when "10100101110010",
                             4712 when "10100101110011",
                             4712 when "10100101110100",
                             4711 when "10100101110101",
                             4711 when "10100101110110",
                             4710 when "10100101110111",
                             4710 when "10100101111000",
                             4709 when "10100101111001",
                             4709 when "10100101111010",
                             4709 when "10100101111011",
                             4708 when "10100101111100",
                             4708 when "10100101111101",
                             4707 when "10100101111110",
                             4707 when "10100101111111",
                             4706 when "10100110000000",
                             4706 when "10100110000001",
                             4705 when "10100110000010",
                             4705 when "10100110000011",
                             4705 when "10100110000100",
                             4704 when "10100110000101",
                             4704 when "10100110000110",
                             4703 when "10100110000111",
                             4703 when "10100110001000",
                             4702 when "10100110001001",
                             4702 when "10100110001010",
                             4701 when "10100110001011",
                             4701 when "10100110001100",
                             4701 when "10100110001101",
                             4700 when "10100110001110",
                             4700 when "10100110001111",
                             4699 when "10100110010000",
                             4699 when "10100110010001",
                             4698 when "10100110010010",
                             4698 when "10100110010011",
                             4697 when "10100110010100",
                             4697 when "10100110010101",
                             4697 when "10100110010110",
                             4696 when "10100110010111",
                             4696 when "10100110011000",
                             4695 when "10100110011001",
                             4695 when "10100110011010",
                             4694 when "10100110011011",
                             4694 when "10100110011100",
                             4694 when "10100110011101",
                             4693 when "10100110011110",
                             4693 when "10100110011111",
                             4692 when "10100110100000",
                             4692 when "10100110100001",
                             4691 when "10100110100010",
                             4691 when "10100110100011",
                             4690 when "10100110100100",
                             4690 when "10100110100101",
                             4690 when "10100110100110",
                             4689 when "10100110100111",
                             4689 when "10100110101000",
                             4688 when "10100110101001",
                             4688 when "10100110101010",
                             4687 when "10100110101011",
                             4687 when "10100110101100",
                             4686 when "10100110101101",
                             4686 when "10100110101110",
                             4686 when "10100110101111",
                             4685 when "10100110110000",
                             4685 when "10100110110001",
                             4684 when "10100110110010",
                             4684 when "10100110110011",
                             4683 when "10100110110100",
                             4683 when "10100110110101",
                             4683 when "10100110110110",
                             4682 when "10100110110111",
                             4682 when "10100110111000",
                             4681 when "10100110111001",
                             4681 when "10100110111010",
                             4680 when "10100110111011",
                             4680 when "10100110111100",
                             4679 when "10100110111101",
                             4679 when "10100110111110",
                             4679 when "10100110111111",
                             4678 when "10100111000000",
                             4678 when "10100111000001",
                             4677 when "10100111000010",
                             4677 when "10100111000011",
                             4676 when "10100111000100",
                             4676 when "10100111000101",
                             4676 when "10100111000110",
                             4675 when "10100111000111",
                             4675 when "10100111001000",
                             4674 when "10100111001001",
                             4674 when "10100111001010",
                             4673 when "10100111001011",
                             4673 when "10100111001100",
                             4672 when "10100111001101",
                             4672 when "10100111001110",
                             4672 when "10100111001111",
                             4671 when "10100111010000",
                             4671 when "10100111010001",
                             4670 when "10100111010010",
                             4670 when "10100111010011",
                             4669 when "10100111010100",
                             4669 when "10100111010101",
                             4669 when "10100111010110",
                             4668 when "10100111010111",
                             4668 when "10100111011000",
                             4667 when "10100111011001",
                             4667 when "10100111011010",
                             4666 when "10100111011011",
                             4666 when "10100111011100",
                             4665 when "10100111011101",
                             4665 when "10100111011110",
                             4665 when "10100111011111",
                             4664 when "10100111100000",
                             4664 when "10100111100001",
                             4663 when "10100111100010",
                             4663 when "10100111100011",
                             4662 when "10100111100100",
                             4662 when "10100111100101",
                             4662 when "10100111100110",
                             4661 when "10100111100111",
                             4661 when "10100111101000",
                             4660 when "10100111101001",
                             4660 when "10100111101010",
                             4659 when "10100111101011",
                             4659 when "10100111101100",
                             4659 when "10100111101101",
                             4658 when "10100111101110",
                             4658 when "10100111101111",
                             4657 when "10100111110000",
                             4657 when "10100111110001",
                             4656 when "10100111110010",
                             4656 when "10100111110011",
                             4655 when "10100111110100",
                             4655 when "10100111110101",
                             4655 when "10100111110110",
                             4654 when "10100111110111",
                             4654 when "10100111111000",
                             4653 when "10100111111001",
                             4653 when "10100111111010",
                             4652 when "10100111111011",
                             4652 when "10100111111100",
                             4652 when "10100111111101",
                             4651 when "10100111111110",
                             4651 when "10100111111111",
                             4650 when "10101000000000",
                             4650 when "10101000000001",
                             4649 when "10101000000010",
                             4649 when "10101000000011",
                             4649 when "10101000000100",
                             4648 when "10101000000101",
                             4648 when "10101000000110",
                             4647 when "10101000000111",
                             4647 when "10101000001000",
                             4646 when "10101000001001",
                             4646 when "10101000001010",
                             4646 when "10101000001011",
                             4645 when "10101000001100",
                             4645 when "10101000001101",
                             4644 when "10101000001110",
                             4644 when "10101000001111",
                             4643 when "10101000010000",
                             4643 when "10101000010001",
                             4643 when "10101000010010",
                             4642 when "10101000010011",
                             4642 when "10101000010100",
                             4641 when "10101000010101",
                             4641 when "10101000010110",
                             4640 when "10101000010111",
                             4640 when "10101000011000",
                             4640 when "10101000011001",
                             4639 when "10101000011010",
                             4639 when "10101000011011",
                             4638 when "10101000011100",
                             4638 when "10101000011101",
                             4637 when "10101000011110",
                             4637 when "10101000011111",
                             4636 when "10101000100000",
                             4636 when "10101000100001",
                             4636 when "10101000100010",
                             4635 when "10101000100011",
                             4635 when "10101000100100",
                             4634 when "10101000100101",
                             4634 when "10101000100110",
                             4633 when "10101000100111",
                             4633 when "10101000101000",
                             4633 when "10101000101001",
                             4632 when "10101000101010",
                             4632 when "10101000101011",
                             4631 when "10101000101100",
                             4631 when "10101000101101",
                             4630 when "10101000101110",
                             4630 when "10101000101111",
                             4630 when "10101000110000",
                             4629 when "10101000110001",
                             4629 when "10101000110010",
                             4628 when "10101000110011",
                             4628 when "10101000110100",
                             4627 when "10101000110101",
                             4627 when "10101000110110",
                             4627 when "10101000110111",
                             4626 when "10101000111000",
                             4626 when "10101000111001",
                             4625 when "10101000111010",
                             4625 when "10101000111011",
                             4624 when "10101000111100",
                             4624 when "10101000111101",
                             4624 when "10101000111110",
                             4623 when "10101000111111",
                             4623 when "10101001000000",
                             4622 when "10101001000001",
                             4622 when "10101001000010",
                             4621 when "10101001000011",
                             4621 when "10101001000100",
                             4621 when "10101001000101",
                             4620 when "10101001000110",
                             4620 when "10101001000111",
                             4619 when "10101001001000",
                             4619 when "10101001001001",
                             4619 when "10101001001010",
                             4618 when "10101001001011",
                             4618 when "10101001001100",
                             4617 when "10101001001101",
                             4617 when "10101001001110",
                             4616 when "10101001001111",
                             4616 when "10101001010000",
                             4616 when "10101001010001",
                             4615 when "10101001010010",
                             4615 when "10101001010011",
                             4614 when "10101001010100",
                             4614 when "10101001010101",
                             4613 when "10101001010110",
                             4613 when "10101001010111",
                             4613 when "10101001011000",
                             4612 when "10101001011001",
                             4612 when "10101001011010",
                             4611 when "10101001011011",
                             4611 when "10101001011100",
                             4610 when "10101001011101",
                             4610 when "10101001011110",
                             4610 when "10101001011111",
                             4609 when "10101001100000",
                             4609 when "10101001100001",
                             4608 when "10101001100010",
                             4608 when "10101001100011",
                             4607 when "10101001100100",
                             4607 when "10101001100101",
                             4607 when "10101001100110",
                             4606 when "10101001100111",
                             4606 when "10101001101000",
                             4605 when "10101001101001",
                             4605 when "10101001101010",
                             4604 when "10101001101011",
                             4604 when "10101001101100",
                             4604 when "10101001101101",
                             4603 when "10101001101110",
                             4603 when "10101001101111",
                             4602 when "10101001110000",
                             4602 when "10101001110001",
                             4602 when "10101001110010",
                             4601 when "10101001110011",
                             4601 when "10101001110100",
                             4600 when "10101001110101",
                             4600 when "10101001110110",
                             4599 when "10101001110111",
                             4599 when "10101001111000",
                             4599 when "10101001111001",
                             4598 when "10101001111010",
                             4598 when "10101001111011",
                             4597 when "10101001111100",
                             4597 when "10101001111101",
                             4596 when "10101001111110",
                             4596 when "10101001111111",
                             4596 when "10101010000000",
                             4595 when "10101010000001",
                             4595 when "10101010000010",
                             4594 when "10101010000011",
                             4594 when "10101010000100",
                             4593 when "10101010000101",
                             4593 when "10101010000110",
                             4593 when "10101010000111",
                             4592 when "10101010001000",
                             4592 when "10101010001001",
                             4591 when "10101010001010",
                             4591 when "10101010001011",
                             4591 when "10101010001100",
                             4590 when "10101010001101",
                             4590 when "10101010001110",
                             4589 when "10101010001111",
                             4589 when "10101010010000",
                             4588 when "10101010010001",
                             4588 when "10101010010010",
                             4588 when "10101010010011",
                             4587 when "10101010010100",
                             4587 when "10101010010101",
                             4586 when "10101010010110",
                             4586 when "10101010010111",
                             4585 when "10101010011000",
                             4585 when "10101010011001",
                             4585 when "10101010011010",
                             4584 when "10101010011011",
                             4584 when "10101010011100",
                             4583 when "10101010011101",
                             4583 when "10101010011110",
                             4583 when "10101010011111",
                             4582 when "10101010100000",
                             4582 when "10101010100001",
                             4581 when "10101010100010",
                             4581 when "10101010100011",
                             4580 when "10101010100100",
                             4580 when "10101010100101",
                             4580 when "10101010100110",
                             4579 when "10101010100111",
                             4579 when "10101010101000",
                             4578 when "10101010101001",
                             4578 when "10101010101010",
                             4577 when "10101010101011",
                             4577 when "10101010101100",
                             4577 when "10101010101101",
                             4576 when "10101010101110",
                             4576 when "10101010101111",
                             4575 when "10101010110000",
                             4575 when "10101010110001",
                             4575 when "10101010110010",
                             4574 when "10101010110011",
                             4574 when "10101010110100",
                             4573 when "10101010110101",
                             4573 when "10101010110110",
                             4572 when "10101010110111",
                             4572 when "10101010111000",
                             4572 when "10101010111001",
                             4571 when "10101010111010",
                             4571 when "10101010111011",
                             4570 when "10101010111100",
                             4570 when "10101010111101",
                             4570 when "10101010111110",
                             4569 when "10101010111111",
                             4569 when "10101011000000",
                             4568 when "10101011000001",
                             4568 when "10101011000010",
                             4567 when "10101011000011",
                             4567 when "10101011000100",
                             4567 when "10101011000101",
                             4566 when "10101011000110",
                             4566 when "10101011000111",
                             4565 when "10101011001000",
                             4565 when "10101011001001",
                             4565 when "10101011001010",
                             4564 when "10101011001011",
                             4564 when "10101011001100",
                             4563 when "10101011001101",
                             4563 when "10101011001110",
                             4562 when "10101011001111",
                             4562 when "10101011010000",
                             4562 when "10101011010001",
                             4561 when "10101011010010",
                             4561 when "10101011010011",
                             4560 when "10101011010100",
                             4560 when "10101011010101",
                             4560 when "10101011010110",
                             4559 when "10101011010111",
                             4559 when "10101011011000",
                             4558 when "10101011011001",
                             4558 when "10101011011010",
                             4557 when "10101011011011",
                             4557 when "10101011011100",
                             4557 when "10101011011101",
                             4556 when "10101011011110",
                             4556 when "10101011011111",
                             4555 when "10101011100000",
                             4555 when "10101011100001",
                             4555 when "10101011100010",
                             4554 when "10101011100011",
                             4554 when "10101011100100",
                             4553 when "10101011100101",
                             4553 when "10101011100110",
                             4552 when "10101011100111",
                             4552 when "10101011101000",
                             4552 when "10101011101001",
                             4551 when "10101011101010",
                             4551 when "10101011101011",
                             4550 when "10101011101100",
                             4550 when "10101011101101",
                             4550 when "10101011101110",
                             4549 when "10101011101111",
                             4549 when "10101011110000",
                             4548 when "10101011110001",
                             4548 when "10101011110010",
                             4548 when "10101011110011",
                             4547 when "10101011110100",
                             4547 when "10101011110101",
                             4546 when "10101011110110",
                             4546 when "10101011110111",
                             4545 when "10101011111000",
                             4545 when "10101011111001",
                             4545 when "10101011111010",
                             4544 when "10101011111011",
                             4544 when "10101011111100",
                             4543 when "10101011111101",
                             4543 when "10101011111110",
                             4543 when "10101011111111",
                             4542 when "10101100000000",
                             4542 when "10101100000001",
                             4541 when "10101100000010",
                             4541 when "10101100000011",
                             4541 when "10101100000100",
                             4540 when "10101100000101",
                             4540 when "10101100000110",
                             4539 when "10101100000111",
                             4539 when "10101100001000",
                             4538 when "10101100001001",
                             4538 when "10101100001010",
                             4538 when "10101100001011",
                             4537 when "10101100001100",
                             4537 when "10101100001101",
                             4536 when "10101100001110",
                             4536 when "10101100001111",
                             4536 when "10101100010000",
                             4535 when "10101100010001",
                             4535 when "10101100010010",
                             4534 when "10101100010011",
                             4534 when "10101100010100",
                             4534 when "10101100010101",
                             4533 when "10101100010110",
                             4533 when "10101100010111",
                             4532 when "10101100011000",
                             4532 when "10101100011001",
                             4531 when "10101100011010",
                             4531 when "10101100011011",
                             4531 when "10101100011100",
                             4530 when "10101100011101",
                             4530 when "10101100011110",
                             4529 when "10101100011111",
                             4529 when "10101100100000",
                             4529 when "10101100100001",
                             4528 when "10101100100010",
                             4528 when "10101100100011",
                             4527 when "10101100100100",
                             4527 when "10101100100101",
                             4527 when "10101100100110",
                             4526 when "10101100100111",
                             4526 when "10101100101000",
                             4525 when "10101100101001",
                             4525 when "10101100101010",
                             4524 when "10101100101011",
                             4524 when "10101100101100",
                             4524 when "10101100101101",
                             4523 when "10101100101110",
                             4523 when "10101100101111",
                             4522 when "10101100110000",
                             4522 when "10101100110001",
                             4522 when "10101100110010",
                             4521 when "10101100110011",
                             4521 when "10101100110100",
                             4520 when "10101100110101",
                             4520 when "10101100110110",
                             4520 when "10101100110111",
                             4519 when "10101100111000",
                             4519 when "10101100111001",
                             4518 when "10101100111010",
                             4518 when "10101100111011",
                             4518 when "10101100111100",
                             4517 when "10101100111101",
                             4517 when "10101100111110",
                             4516 when "10101100111111",
                             4516 when "10101101000000",
                             4515 when "10101101000001",
                             4515 when "10101101000010",
                             4515 when "10101101000011",
                             4514 when "10101101000100",
                             4514 when "10101101000101",
                             4513 when "10101101000110",
                             4513 when "10101101000111",
                             4513 when "10101101001000",
                             4512 when "10101101001001",
                             4512 when "10101101001010",
                             4511 when "10101101001011",
                             4511 when "10101101001100",
                             4511 when "10101101001101",
                             4510 when "10101101001110",
                             4510 when "10101101001111",
                             4509 when "10101101010000",
                             4509 when "10101101010001",
                             4509 when "10101101010010",
                             4508 when "10101101010011",
                             4508 when "10101101010100",
                             4507 when "10101101010101",
                             4507 when "10101101010110",
                             4507 when "10101101010111",
                             4506 when "10101101011000",
                             4506 when "10101101011001",
                             4505 when "10101101011010",
                             4505 when "10101101011011",
                             4505 when "10101101011100",
                             4504 when "10101101011101",
                             4504 when "10101101011110",
                             4503 when "10101101011111",
                             4503 when "10101101100000",
                             4502 when "10101101100001",
                             4502 when "10101101100010",
                             4502 when "10101101100011",
                             4501 when "10101101100100",
                             4501 when "10101101100101",
                             4500 when "10101101100110",
                             4500 when "10101101100111",
                             4500 when "10101101101000",
                             4499 when "10101101101001",
                             4499 when "10101101101010",
                             4498 when "10101101101011",
                             4498 when "10101101101100",
                             4498 when "10101101101101",
                             4497 when "10101101101110",
                             4497 when "10101101101111",
                             4496 when "10101101110000",
                             4496 when "10101101110001",
                             4496 when "10101101110010",
                             4495 when "10101101110011",
                             4495 when "10101101110100",
                             4494 when "10101101110101",
                             4494 when "10101101110110",
                             4494 when "10101101110111",
                             4493 when "10101101111000",
                             4493 when "10101101111001",
                             4492 when "10101101111010",
                             4492 when "10101101111011",
                             4492 when "10101101111100",
                             4491 when "10101101111101",
                             4491 when "10101101111110",
                             4490 when "10101101111111",
                             4490 when "10101110000000",
                             4490 when "10101110000001",
                             4489 when "10101110000010",
                             4489 when "10101110000011",
                             4488 when "10101110000100",
                             4488 when "10101110000101",
                             4488 when "10101110000110",
                             4487 when "10101110000111",
                             4487 when "10101110001000",
                             4486 when "10101110001001",
                             4486 when "10101110001010",
                             4486 when "10101110001011",
                             4485 when "10101110001100",
                             4485 when "10101110001101",
                             4484 when "10101110001110",
                             4484 when "10101110001111",
                             4484 when "10101110010000",
                             4483 when "10101110010001",
                             4483 when "10101110010010",
                             4482 when "10101110010011",
                             4482 when "10101110010100",
                             4481 when "10101110010101",
                             4481 when "10101110010110",
                             4481 when "10101110010111",
                             4480 when "10101110011000",
                             4480 when "10101110011001",
                             4479 when "10101110011010",
                             4479 when "10101110011011",
                             4479 when "10101110011100",
                             4478 when "10101110011101",
                             4478 when "10101110011110",
                             4477 when "10101110011111",
                             4477 when "10101110100000",
                             4477 when "10101110100001",
                             4476 when "10101110100010",
                             4476 when "10101110100011",
                             4475 when "10101110100100",
                             4475 when "10101110100101",
                             4475 when "10101110100110",
                             4474 when "10101110100111",
                             4474 when "10101110101000",
                             4473 when "10101110101001",
                             4473 when "10101110101010",
                             4473 when "10101110101011",
                             4472 when "10101110101100",
                             4472 when "10101110101101",
                             4471 when "10101110101110",
                             4471 when "10101110101111",
                             4471 when "10101110110000",
                             4470 when "10101110110001",
                             4470 when "10101110110010",
                             4469 when "10101110110011",
                             4469 when "10101110110100",
                             4469 when "10101110110101",
                             4468 when "10101110110110",
                             4468 when "10101110110111",
                             4467 when "10101110111000",
                             4467 when "10101110111001",
                             4467 when "10101110111010",
                             4466 when "10101110111011",
                             4466 when "10101110111100",
                             4465 when "10101110111101",
                             4465 when "10101110111110",
                             4465 when "10101110111111",
                             4464 when "10101111000000",
                             4464 when "10101111000001",
                             4463 when "10101111000010",
                             4463 when "10101111000011",
                             4463 when "10101111000100",
                             4462 when "10101111000101",
                             4462 when "10101111000110",
                             4461 when "10101111000111",
                             4461 when "10101111001000",
                             4461 when "10101111001001",
                             4460 when "10101111001010",
                             4460 when "10101111001011",
                             4460 when "10101111001100",
                             4459 when "10101111001101",
                             4459 when "10101111001110",
                             4458 when "10101111001111",
                             4458 when "10101111010000",
                             4458 when "10101111010001",
                             4457 when "10101111010010",
                             4457 when "10101111010011",
                             4456 when "10101111010100",
                             4456 when "10101111010101",
                             4456 when "10101111010110",
                             4455 when "10101111010111",
                             4455 when "10101111011000",
                             4454 when "10101111011001",
                             4454 when "10101111011010",
                             4454 when "10101111011011",
                             4453 when "10101111011100",
                             4453 when "10101111011101",
                             4452 when "10101111011110",
                             4452 when "10101111011111",
                             4452 when "10101111100000",
                             4451 when "10101111100001",
                             4451 when "10101111100010",
                             4450 when "10101111100011",
                             4450 when "10101111100100",
                             4450 when "10101111100101",
                             4449 when "10101111100110",
                             4449 when "10101111100111",
                             4448 when "10101111101000",
                             4448 when "10101111101001",
                             4448 when "10101111101010",
                             4447 when "10101111101011",
                             4447 when "10101111101100",
                             4446 when "10101111101101",
                             4446 when "10101111101110",
                             4446 when "10101111101111",
                             4445 when "10101111110000",
                             4445 when "10101111110001",
                             4444 when "10101111110010",
                             4444 when "10101111110011",
                             4444 when "10101111110100",
                             4443 when "10101111110101",
                             4443 when "10101111110110",
                             4442 when "10101111110111",
                             4442 when "10101111111000",
                             4442 when "10101111111001",
                             4441 when "10101111111010",
                             4441 when "10101111111011",
                             4440 when "10101111111100",
                             4440 when "10101111111101",
                             4440 when "10101111111110",
                             4439 when "10101111111111",
                             4439 when "10110000000000",
                             4439 when "10110000000001",
                             4438 when "10110000000010",
                             4438 when "10110000000011",
                             4437 when "10110000000100",
                             4437 when "10110000000101",
                             4437 when "10110000000110",
                             4436 when "10110000000111",
                             4436 when "10110000001000",
                             4435 when "10110000001001",
                             4435 when "10110000001010",
                             4435 when "10110000001011",
                             4434 when "10110000001100",
                             4434 when "10110000001101",
                             4433 when "10110000001110",
                             4433 when "10110000001111",
                             4433 when "10110000010000",
                             4432 when "10110000010001",
                             4432 when "10110000010010",
                             4431 when "10110000010011",
                             4431 when "10110000010100",
                             4431 when "10110000010101",
                             4430 when "10110000010110",
                             4430 when "10110000010111",
                             4429 when "10110000011000",
                             4429 when "10110000011001",
                             4429 when "10110000011010",
                             4428 when "10110000011011",
                             4428 when "10110000011100",
                             4428 when "10110000011101",
                             4427 when "10110000011110",
                             4427 when "10110000011111",
                             4426 when "10110000100000",
                             4426 when "10110000100001",
                             4426 when "10110000100010",
                             4425 when "10110000100011",
                             4425 when "10110000100100",
                             4424 when "10110000100101",
                             4424 when "10110000100110",
                             4424 when "10110000100111",
                             4423 when "10110000101000",
                             4423 when "10110000101001",
                             4422 when "10110000101010",
                             4422 when "10110000101011",
                             4422 when "10110000101100",
                             4421 when "10110000101101",
                             4421 when "10110000101110",
                             4420 when "10110000101111",
                             4420 when "10110000110000",
                             4420 when "10110000110001",
                             4419 when "10110000110010",
                             4419 when "10110000110011",
                             4419 when "10110000110100",
                             4418 when "10110000110101",
                             4418 when "10110000110110",
                             4417 when "10110000110111",
                             4417 when "10110000111000",
                             4417 when "10110000111001",
                             4416 when "10110000111010",
                             4416 when "10110000111011",
                             4415 when "10110000111100",
                             4415 when "10110000111101",
                             4415 when "10110000111110",
                             4414 when "10110000111111",
                             4414 when "10110001000000",
                             4413 when "10110001000001",
                             4413 when "10110001000010",
                             4413 when "10110001000011",
                             4412 when "10110001000100",
                             4412 when "10110001000101",
                             4412 when "10110001000110",
                             4411 when "10110001000111",
                             4411 when "10110001001000",
                             4410 when "10110001001001",
                             4410 when "10110001001010",
                             4410 when "10110001001011",
                             4409 when "10110001001100",
                             4409 when "10110001001101",
                             4408 when "10110001001110",
                             4408 when "10110001001111",
                             4408 when "10110001010000",
                             4407 when "10110001010001",
                             4407 when "10110001010010",
                             4406 when "10110001010011",
                             4406 when "10110001010100",
                             4406 when "10110001010101",
                             4405 when "10110001010110",
                             4405 when "10110001010111",
                             4405 when "10110001011000",
                             4404 when "10110001011001",
                             4404 when "10110001011010",
                             4403 when "10110001011011",
                             4403 when "10110001011100",
                             4403 when "10110001011101",
                             4402 when "10110001011110",
                             4402 when "10110001011111",
                             4401 when "10110001100000",
                             4401 when "10110001100001",
                             4401 when "10110001100010",
                             4400 when "10110001100011",
                             4400 when "10110001100100",
                             4399 when "10110001100101",
                             4399 when "10110001100110",
                             4399 when "10110001100111",
                             4398 when "10110001101000",
                             4398 when "10110001101001",
                             4398 when "10110001101010",
                             4397 when "10110001101011",
                             4397 when "10110001101100",
                             4396 when "10110001101101",
                             4396 when "10110001101110",
                             4396 when "10110001101111",
                             4395 when "10110001110000",
                             4395 when "10110001110001",
                             4394 when "10110001110010",
                             4394 when "10110001110011",
                             4394 when "10110001110100",
                             4393 when "10110001110101",
                             4393 when "10110001110110",
                             4393 when "10110001110111",
                             4392 when "10110001111000",
                             4392 when "10110001111001",
                             4391 when "10110001111010",
                             4391 when "10110001111011",
                             4391 when "10110001111100",
                             4390 when "10110001111101",
                             4390 when "10110001111110",
                             4389 when "10110001111111",
                             4389 when "10110010000000",
                             4389 when "10110010000001",
                             4388 when "10110010000010",
                             4388 when "10110010000011",
                             4388 when "10110010000100",
                             4387 when "10110010000101",
                             4387 when "10110010000110",
                             4386 when "10110010000111",
                             4386 when "10110010001000",
                             4386 when "10110010001001",
                             4385 when "10110010001010",
                             4385 when "10110010001011",
                             4384 when "10110010001100",
                             4384 when "10110010001101",
                             4384 when "10110010001110",
                             4383 when "10110010001111",
                             4383 when "10110010010000",
                             4383 when "10110010010001",
                             4382 when "10110010010010",
                             4382 when "10110010010011",
                             4381 when "10110010010100",
                             4381 when "10110010010101",
                             4381 when "10110010010110",
                             4380 when "10110010010111",
                             4380 when "10110010011000",
                             4379 when "10110010011001",
                             4379 when "10110010011010",
                             4379 when "10110010011011",
                             4378 when "10110010011100",
                             4378 when "10110010011101",
                             4378 when "10110010011110",
                             4377 when "10110010011111",
                             4377 when "10110010100000",
                             4376 when "10110010100001",
                             4376 when "10110010100010",
                             4376 when "10110010100011",
                             4375 when "10110010100100",
                             4375 when "10110010100101",
                             4374 when "10110010100110",
                             4374 when "10110010100111",
                             4374 when "10110010101000",
                             4373 when "10110010101001",
                             4373 when "10110010101010",
                             4373 when "10110010101011",
                             4372 when "10110010101100",
                             4372 when "10110010101101",
                             4371 when "10110010101110",
                             4371 when "10110010101111",
                             4371 when "10110010110000",
                             4370 when "10110010110001",
                             4370 when "10110010110010",
                             4369 when "10110010110011",
                             4369 when "10110010110100",
                             4369 when "10110010110101",
                             4368 when "10110010110110",
                             4368 when "10110010110111",
                             4368 when "10110010111000",
                             4367 when "10110010111001",
                             4367 when "10110010111010",
                             4366 when "10110010111011",
                             4366 when "10110010111100",
                             4366 when "10110010111101",
                             4365 when "10110010111110",
                             4365 when "10110010111111",
                             4365 when "10110011000000",
                             4364 when "10110011000001",
                             4364 when "10110011000010",
                             4363 when "10110011000011",
                             4363 when "10110011000100",
                             4363 when "10110011000101",
                             4362 when "10110011000110",
                             4362 when "10110011000111",
                             4361 when "10110011001000",
                             4361 when "10110011001001",
                             4361 when "10110011001010",
                             4360 when "10110011001011",
                             4360 when "10110011001100",
                             4360 when "10110011001101",
                             4359 when "10110011001110",
                             4359 when "10110011001111",
                             4358 when "10110011010000",
                             4358 when "10110011010001",
                             4358 when "10110011010010",
                             4357 when "10110011010011",
                             4357 when "10110011010100",
                             4357 when "10110011010101",
                             4356 when "10110011010110",
                             4356 when "10110011010111",
                             4355 when "10110011011000",
                             4355 when "10110011011001",
                             4355 when "10110011011010",
                             4354 when "10110011011011",
                             4354 when "10110011011100",
                             4354 when "10110011011101",
                             4353 when "10110011011110",
                             4353 when "10110011011111",
                             4352 when "10110011100000",
                             4352 when "10110011100001",
                             4352 when "10110011100010",
                             4351 when "10110011100011",
                             4351 when "10110011100100",
                             4350 when "10110011100101",
                             4350 when "10110011100110",
                             4350 when "10110011100111",
                             4349 when "10110011101000",
                             4349 when "10110011101001",
                             4349 when "10110011101010",
                             4348 when "10110011101011",
                             4348 when "10110011101100",
                             4347 when "10110011101101",
                             4347 when "10110011101110",
                             4347 when "10110011101111",
                             4346 when "10110011110000",
                             4346 when "10110011110001",
                             4346 when "10110011110010",
                             4345 when "10110011110011",
                             4345 when "10110011110100",
                             4344 when "10110011110101",
                             4344 when "10110011110110",
                             4344 when "10110011110111",
                             4343 when "10110011111000",
                             4343 when "10110011111001",
                             4343 when "10110011111010",
                             4342 when "10110011111011",
                             4342 when "10110011111100",
                             4341 when "10110011111101",
                             4341 when "10110011111110",
                             4341 when "10110011111111",
                             4340 when "10110100000000",
                             4340 when "10110100000001",
                             4340 when "10110100000010",
                             4339 when "10110100000011",
                             4339 when "10110100000100",
                             4338 when "10110100000101",
                             4338 when "10110100000110",
                             4338 when "10110100000111",
                             4337 when "10110100001000",
                             4337 when "10110100001001",
                             4337 when "10110100001010",
                             4336 when "10110100001011",
                             4336 when "10110100001100",
                             4335 when "10110100001101",
                             4335 when "10110100001110",
                             4335 when "10110100001111",
                             4334 when "10110100010000",
                             4334 when "10110100010001",
                             4334 when "10110100010010",
                             4333 when "10110100010011",
                             4333 when "10110100010100",
                             4332 when "10110100010101",
                             4332 when "10110100010110",
                             4332 when "10110100010111",
                             4331 when "10110100011000",
                             4331 when "10110100011001",
                             4331 when "10110100011010",
                             4330 when "10110100011011",
                             4330 when "10110100011100",
                             4329 when "10110100011101",
                             4329 when "10110100011110",
                             4329 when "10110100011111",
                             4328 when "10110100100000",
                             4328 when "10110100100001",
                             4328 when "10110100100010",
                             4327 when "10110100100011",
                             4327 when "10110100100100",
                             4326 when "10110100100101",
                             4326 when "10110100100110",
                             4326 when "10110100100111",
                             4325 when "10110100101000",
                             4325 when "10110100101001",
                             4325 when "10110100101010",
                             4324 when "10110100101011",
                             4324 when "10110100101100",
                             4323 when "10110100101101",
                             4323 when "10110100101110",
                             4323 when "10110100101111",
                             4322 when "10110100110000",
                             4322 when "10110100110001",
                             4322 when "10110100110010",
                             4321 when "10110100110011",
                             4321 when "10110100110100",
                             4320 when "10110100110101",
                             4320 when "10110100110110",
                             4320 when "10110100110111",
                             4319 when "10110100111000",
                             4319 when "10110100111001",
                             4319 when "10110100111010",
                             4318 when "10110100111011",
                             4318 when "10110100111100",
                             4317 when "10110100111101",
                             4317 when "10110100111110",
                             4317 when "10110100111111",
                             4316 when "10110101000000",
                             4316 when "10110101000001",
                             4316 when "10110101000010",
                             4315 when "10110101000011",
                             4315 when "10110101000100",
                             4314 when "10110101000101",
                             4314 when "10110101000110",
                             4314 when "10110101000111",
                             4313 when "10110101001000",
                             4313 when "10110101001001",
                             4313 when "10110101001010",
                             4312 when "10110101001011",
                             4312 when "10110101001100",
                             4311 when "10110101001101",
                             4311 when "10110101001110",
                             4311 when "10110101001111",
                             4310 when "10110101010000",
                             4310 when "10110101010001",
                             4310 when "10110101010010",
                             4309 when "10110101010011",
                             4309 when "10110101010100",
                             4308 when "10110101010101",
                             4308 when "10110101010110",
                             4308 when "10110101010111",
                             4307 when "10110101011000",
                             4307 when "10110101011001",
                             4307 when "10110101011010",
                             4306 when "10110101011011",
                             4306 when "10110101011100",
                             4306 when "10110101011101",
                             4305 when "10110101011110",
                             4305 when "10110101011111",
                             4304 when "10110101100000",
                             4304 when "10110101100001",
                             4304 when "10110101100010",
                             4303 when "10110101100011",
                             4303 when "10110101100100",
                             4303 when "10110101100101",
                             4302 when "10110101100110",
                             4302 when "10110101100111",
                             4301 when "10110101101000",
                             4301 when "10110101101001",
                             4301 when "10110101101010",
                             4300 when "10110101101011",
                             4300 when "10110101101100",
                             4300 when "10110101101101",
                             4299 when "10110101101110",
                             4299 when "10110101101111",
                             4298 when "10110101110000",
                             4298 when "10110101110001",
                             4298 when "10110101110010",
                             4297 when "10110101110011",
                             4297 when "10110101110100",
                             4297 when "10110101110101",
                             4296 when "10110101110110",
                             4296 when "10110101110111",
                             4296 when "10110101111000",
                             4295 when "10110101111001",
                             4295 when "10110101111010",
                             4294 when "10110101111011",
                             4294 when "10110101111100",
                             4294 when "10110101111101",
                             4293 when "10110101111110",
                             4293 when "10110101111111",
                             4293 when "10110110000000",
                             4292 when "10110110000001",
                             4292 when "10110110000010",
                             4291 when "10110110000011",
                             4291 when "10110110000100",
                             4291 when "10110110000101",
                             4290 when "10110110000110",
                             4290 when "10110110000111",
                             4290 when "10110110001000",
                             4289 when "10110110001001",
                             4289 when "10110110001010",
                             4289 when "10110110001011",
                             4288 when "10110110001100",
                             4288 when "10110110001101",
                             4287 when "10110110001110",
                             4287 when "10110110001111",
                             4287 when "10110110010000",
                             4286 when "10110110010001",
                             4286 when "10110110010010",
                             4286 when "10110110010011",
                             4285 when "10110110010100",
                             4285 when "10110110010101",
                             4284 when "10110110010110",
                             4284 when "10110110010111",
                             4284 when "10110110011000",
                             4283 when "10110110011001",
                             4283 when "10110110011010",
                             4283 when "10110110011011",
                             4282 when "10110110011100",
                             4282 when "10110110011101",
                             4282 when "10110110011110",
                             4281 when "10110110011111",
                             4281 when "10110110100000",
                             4280 when "10110110100001",
                             4280 when "10110110100010",
                             4280 when "10110110100011",
                             4279 when "10110110100100",
                             4279 when "10110110100101",
                             4279 when "10110110100110",
                             4278 when "10110110100111",
                             4278 when "10110110101000",
                             4278 when "10110110101001",
                             4277 when "10110110101010",
                             4277 when "10110110101011",
                             4276 when "10110110101100",
                             4276 when "10110110101101",
                             4276 when "10110110101110",
                             4275 when "10110110101111",
                             4275 when "10110110110000",
                             4275 when "10110110110001",
                             4274 when "10110110110010",
                             4274 when "10110110110011",
                             4274 when "10110110110100",
                             4273 when "10110110110101",
                             4273 when "10110110110110",
                             4272 when "10110110110111",
                             4272 when "10110110111000",
                             4272 when "10110110111001",
                             4271 when "10110110111010",
                             4271 when "10110110111011",
                             4271 when "10110110111100",
                             4270 when "10110110111101",
                             4270 when "10110110111110",
                             4269 when "10110110111111",
                             4269 when "10110111000000",
                             4269 when "10110111000001",
                             4268 when "10110111000010",
                             4268 when "10110111000011",
                             4268 when "10110111000100",
                             4267 when "10110111000101",
                             4267 when "10110111000110",
                             4267 when "10110111000111",
                             4266 when "10110111001000",
                             4266 when "10110111001001",
                             4265 when "10110111001010",
                             4265 when "10110111001011",
                             4265 when "10110111001100",
                             4264 when "10110111001101",
                             4264 when "10110111001110",
                             4264 when "10110111001111",
                             4263 when "10110111010000",
                             4263 when "10110111010001",
                             4263 when "10110111010010",
                             4262 when "10110111010011",
                             4262 when "10110111010100",
                             4261 when "10110111010101",
                             4261 when "10110111010110",
                             4261 when "10110111010111",
                             4260 when "10110111011000",
                             4260 when "10110111011001",
                             4260 when "10110111011010",
                             4259 when "10110111011011",
                             4259 when "10110111011100",
                             4259 when "10110111011101",
                             4258 when "10110111011110",
                             4258 when "10110111011111",
                             4257 when "10110111100000",
                             4257 when "10110111100001",
                             4257 when "10110111100010",
                             4256 when "10110111100011",
                             4256 when "10110111100100",
                             4256 when "10110111100101",
                             4255 when "10110111100110",
                             4255 when "10110111100111",
                             4255 when "10110111101000",
                             4254 when "10110111101001",
                             4254 when "10110111101010",
                             4254 when "10110111101011",
                             4253 when "10110111101100",
                             4253 when "10110111101101",
                             4252 when "10110111101110",
                             4252 when "10110111101111",
                             4252 when "10110111110000",
                             4251 when "10110111110001",
                             4251 when "10110111110010",
                             4251 when "10110111110011",
                             4250 when "10110111110100",
                             4250 when "10110111110101",
                             4250 when "10110111110110",
                             4249 when "10110111110111",
                             4249 when "10110111111000",
                             4248 when "10110111111001",
                             4248 when "10110111111010",
                             4248 when "10110111111011",
                             4247 when "10110111111100",
                             4247 when "10110111111101",
                             4247 when "10110111111110",
                             4246 when "10110111111111",
                             4246 when "10111000000000",
                             4246 when "10111000000001",
                             4245 when "10111000000010",
                             4245 when "10111000000011",
                             4244 when "10111000000100",
                             4244 when "10111000000101",
                             4244 when "10111000000110",
                             4243 when "10111000000111",
                             4243 when "10111000001000",
                             4243 when "10111000001001",
                             4242 when "10111000001010",
                             4242 when "10111000001011",
                             4242 when "10111000001100",
                             4241 when "10111000001101",
                             4241 when "10111000001110",
                             4241 when "10111000001111",
                             4240 when "10111000010000",
                             4240 when "10111000010001",
                             4239 when "10111000010010",
                             4239 when "10111000010011",
                             4239 when "10111000010100",
                             4238 when "10111000010101",
                             4238 when "10111000010110",
                             4238 when "10111000010111",
                             4237 when "10111000011000",
                             4237 when "10111000011001",
                             4237 when "10111000011010",
                             4236 when "10111000011011",
                             4236 when "10111000011100",
                             4235 when "10111000011101",
                             4235 when "10111000011110",
                             4235 when "10111000011111",
                             4234 when "10111000100000",
                             4234 when "10111000100001",
                             4234 when "10111000100010",
                             4233 when "10111000100011",
                             4233 when "10111000100100",
                             4233 when "10111000100101",
                             4232 when "10111000100110",
                             4232 when "10111000100111",
                             4232 when "10111000101000",
                             4231 when "10111000101001",
                             4231 when "10111000101010",
                             4230 when "10111000101011",
                             4230 when "10111000101100",
                             4230 when "10111000101101",
                             4229 when "10111000101110",
                             4229 when "10111000101111",
                             4229 when "10111000110000",
                             4228 when "10111000110001",
                             4228 when "10111000110010",
                             4228 when "10111000110011",
                             4227 when "10111000110100",
                             4227 when "10111000110101",
                             4227 when "10111000110110",
                             4226 when "10111000110111",
                             4226 when "10111000111000",
                             4225 when "10111000111001",
                             4225 when "10111000111010",
                             4225 when "10111000111011",
                             4224 when "10111000111100",
                             4224 when "10111000111101",
                             4224 when "10111000111110",
                             4223 when "10111000111111",
                             4223 when "10111001000000",
                             4223 when "10111001000001",
                             4222 when "10111001000010",
                             4222 when "10111001000011",
                             4222 when "10111001000100",
                             4221 when "10111001000101",
                             4221 when "10111001000110",
                             4220 when "10111001000111",
                             4220 when "10111001001000",
                             4220 when "10111001001001",
                             4219 when "10111001001010",
                             4219 when "10111001001011",
                             4219 when "10111001001100",
                             4218 when "10111001001101",
                             4218 when "10111001001110",
                             4218 when "10111001001111",
                             4217 when "10111001010000",
                             4217 when "10111001010001",
                             4217 when "10111001010010",
                             4216 when "10111001010011",
                             4216 when "10111001010100",
                             4215 when "10111001010101",
                             4215 when "10111001010110",
                             4215 when "10111001010111",
                             4214 when "10111001011000",
                             4214 when "10111001011001",
                             4214 when "10111001011010",
                             4213 when "10111001011011",
                             4213 when "10111001011100",
                             4213 when "10111001011101",
                             4212 when "10111001011110",
                             4212 when "10111001011111",
                             4212 when "10111001100000",
                             4211 when "10111001100001",
                             4211 when "10111001100010",
                             4211 when "10111001100011",
                             4210 when "10111001100100",
                             4210 when "10111001100101",
                             4209 when "10111001100110",
                             4209 when "10111001100111",
                             4209 when "10111001101000",
                             4208 when "10111001101001",
                             4208 when "10111001101010",
                             4208 when "10111001101011",
                             4207 when "10111001101100",
                             4207 when "10111001101101",
                             4207 when "10111001101110",
                             4206 when "10111001101111",
                             4206 when "10111001110000",
                             4206 when "10111001110001",
                             4205 when "10111001110010",
                             4205 when "10111001110011",
                             4205 when "10111001110100",
                             4204 when "10111001110101",
                             4204 when "10111001110110",
                             4203 when "10111001110111",
                             4203 when "10111001111000",
                             4203 when "10111001111001",
                             4202 when "10111001111010",
                             4202 when "10111001111011",
                             4202 when "10111001111100",
                             4201 when "10111001111101",
                             4201 when "10111001111110",
                             4201 when "10111001111111",
                             4200 when "10111010000000",
                             4200 when "10111010000001",
                             4200 when "10111010000010",
                             4199 when "10111010000011",
                             4199 when "10111010000100",
                             4199 when "10111010000101",
                             4198 when "10111010000110",
                             4198 when "10111010000111",
                             4197 when "10111010001000",
                             4197 when "10111010001001",
                             4197 when "10111010001010",
                             4196 when "10111010001011",
                             4196 when "10111010001100",
                             4196 when "10111010001101",
                             4195 when "10111010001110",
                             4195 when "10111010001111",
                             4195 when "10111010010000",
                             4194 when "10111010010001",
                             4194 when "10111010010010",
                             4194 when "10111010010011",
                             4193 when "10111010010100",
                             4193 when "10111010010101",
                             4193 when "10111010010110",
                             4192 when "10111010010111",
                             4192 when "10111010011000",
                             4191 when "10111010011001",
                             4191 when "10111010011010",
                             4191 when "10111010011011",
                             4190 when "10111010011100",
                             4190 when "10111010011101",
                             4190 when "10111010011110",
                             4189 when "10111010011111",
                             4189 when "10111010100000",
                             4189 when "10111010100001",
                             4188 when "10111010100010",
                             4188 when "10111010100011",
                             4188 when "10111010100100",
                             4187 when "10111010100101",
                             4187 when "10111010100110",
                             4187 when "10111010100111",
                             4186 when "10111010101000",
                             4186 when "10111010101001",
                             4186 when "10111010101010",
                             4185 when "10111010101011",
                             4185 when "10111010101100",
                             4184 when "10111010101101",
                             4184 when "10111010101110",
                             4184 when "10111010101111",
                             4183 when "10111010110000",
                             4183 when "10111010110001",
                             4183 when "10111010110010",
                             4182 when "10111010110011",
                             4182 when "10111010110100",
                             4182 when "10111010110101",
                             4181 when "10111010110110",
                             4181 when "10111010110111",
                             4181 when "10111010111000",
                             4180 when "10111010111001",
                             4180 when "10111010111010",
                             4180 when "10111010111011",
                             4179 when "10111010111100",
                             4179 when "10111010111101",
                             4179 when "10111010111110",
                             4178 when "10111010111111",
                             4178 when "10111011000000",
                             4177 when "10111011000001",
                             4177 when "10111011000010",
                             4177 when "10111011000011",
                             4176 when "10111011000100",
                             4176 when "10111011000101",
                             4176 when "10111011000110",
                             4175 when "10111011000111",
                             4175 when "10111011001000",
                             4175 when "10111011001001",
                             4174 when "10111011001010",
                             4174 when "10111011001011",
                             4174 when "10111011001100",
                             4173 when "10111011001101",
                             4173 when "10111011001110",
                             4173 when "10111011001111",
                             4172 when "10111011010000",
                             4172 when "10111011010001",
                             4172 when "10111011010010",
                             4171 when "10111011010011",
                             4171 when "10111011010100",
                             4170 when "10111011010101",
                             4170 when "10111011010110",
                             4170 when "10111011010111",
                             4169 when "10111011011000",
                             4169 when "10111011011001",
                             4169 when "10111011011010",
                             4168 when "10111011011011",
                             4168 when "10111011011100",
                             4168 when "10111011011101",
                             4167 when "10111011011110",
                             4167 when "10111011011111",
                             4167 when "10111011100000",
                             4166 when "10111011100001",
                             4166 when "10111011100010",
                             4166 when "10111011100011",
                             4165 when "10111011100100",
                             4165 when "10111011100101",
                             4165 when "10111011100110",
                             4164 when "10111011100111",
                             4164 when "10111011101000",
                             4164 when "10111011101001",
                             4163 when "10111011101010",
                             4163 when "10111011101011",
                             4163 when "10111011101100",
                             4162 when "10111011101101",
                             4162 when "10111011101110",
                             4161 when "10111011101111",
                             4161 when "10111011110000",
                             4161 when "10111011110001",
                             4160 when "10111011110010",
                             4160 when "10111011110011",
                             4160 when "10111011110100",
                             4159 when "10111011110101",
                             4159 when "10111011110110",
                             4159 when "10111011110111",
                             4158 when "10111011111000",
                             4158 when "10111011111001",
                             4158 when "10111011111010",
                             4157 when "10111011111011",
                             4157 when "10111011111100",
                             4157 when "10111011111101",
                             4156 when "10111011111110",
                             4156 when "10111011111111",
                             4156 when "10111100000000",
                             4155 when "10111100000001",
                             4155 when "10111100000010",
                             4155 when "10111100000011",
                             4154 when "10111100000100",
                             4154 when "10111100000101",
                             4154 when "10111100000110",
                             4153 when "10111100000111",
                             4153 when "10111100001000",
                             4152 when "10111100001001",
                             4152 when "10111100001010",
                             4152 when "10111100001011",
                             4151 when "10111100001100",
                             4151 when "10111100001101",
                             4151 when "10111100001110",
                             4150 when "10111100001111",
                             4150 when "10111100010000",
                             4150 when "10111100010001",
                             4149 when "10111100010010",
                             4149 when "10111100010011",
                             4149 when "10111100010100",
                             4148 when "10111100010101",
                             4148 when "10111100010110",
                             4148 when "10111100010111",
                             4147 when "10111100011000",
                             4147 when "10111100011001",
                             4147 when "10111100011010",
                             4146 when "10111100011011",
                             4146 when "10111100011100",
                             4146 when "10111100011101",
                             4145 when "10111100011110",
                             4145 when "10111100011111",
                             4145 when "10111100100000",
                             4144 when "10111100100001",
                             4144 when "10111100100010",
                             4144 when "10111100100011",
                             4143 when "10111100100100",
                             4143 when "10111100100101",
                             4143 when "10111100100110",
                             4142 when "10111100100111",
                             4142 when "10111100101000",
                             4141 when "10111100101001",
                             4141 when "10111100101010",
                             4141 when "10111100101011",
                             4140 when "10111100101100",
                             4140 when "10111100101101",
                             4140 when "10111100101110",
                             4139 when "10111100101111",
                             4139 when "10111100110000",
                             4139 when "10111100110001",
                             4138 when "10111100110010",
                             4138 when "10111100110011",
                             4138 when "10111100110100",
                             4137 when "10111100110101",
                             4137 when "10111100110110",
                             4137 when "10111100110111",
                             4136 when "10111100111000",
                             4136 when "10111100111001",
                             4136 when "10111100111010",
                             4135 when "10111100111011",
                             4135 when "10111100111100",
                             4135 when "10111100111101",
                             4134 when "10111100111110",
                             4134 when "10111100111111",
                             4134 when "10111101000000",
                             4133 when "10111101000001",
                             4133 when "10111101000010",
                             4133 when "10111101000011",
                             4132 when "10111101000100",
                             4132 when "10111101000101",
                             4132 when "10111101000110",
                             4131 when "10111101000111",
                             4131 when "10111101001000",
                             4131 when "10111101001001",
                             4130 when "10111101001010",
                             4130 when "10111101001011",
                             4130 when "10111101001100",
                             4129 when "10111101001101",
                             4129 when "10111101001110",
                             4128 when "10111101001111",
                             4128 when "10111101010000",
                             4128 when "10111101010001",
                             4127 when "10111101010010",
                             4127 when "10111101010011",
                             4127 when "10111101010100",
                             4126 when "10111101010101",
                             4126 when "10111101010110",
                             4126 when "10111101010111",
                             4125 when "10111101011000",
                             4125 when "10111101011001",
                             4125 when "10111101011010",
                             4124 when "10111101011011",
                             4124 when "10111101011100",
                             4124 when "10111101011101",
                             4123 when "10111101011110",
                             4123 when "10111101011111",
                             4123 when "10111101100000",
                             4122 when "10111101100001",
                             4122 when "10111101100010",
                             4122 when "10111101100011",
                             4121 when "10111101100100",
                             4121 when "10111101100101",
                             4121 when "10111101100110",
                             4120 when "10111101100111",
                             4120 when "10111101101000",
                             4120 when "10111101101001",
                             4119 when "10111101101010",
                             4119 when "10111101101011",
                             4119 when "10111101101100",
                             4118 when "10111101101101",
                             4118 when "10111101101110",
                             4118 when "10111101101111",
                             4117 when "10111101110000",
                             4117 when "10111101110001",
                             4117 when "10111101110010",
                             4116 when "10111101110011",
                             4116 when "10111101110100",
                             4116 when "10111101110101",
                             4115 when "10111101110110",
                             4115 when "10111101110111",
                             4115 when "10111101111000",
                             4114 when "10111101111001",
                             4114 when "10111101111010",
                             4114 when "10111101111011",
                             4113 when "10111101111100",
                             4113 when "10111101111101",
                             4113 when "10111101111110",
                             4112 when "10111101111111",
                             4112 when "10111110000000",
                             4112 when "10111110000001",
                             4111 when "10111110000010",
                             4111 when "10111110000011",
                             4110 when "10111110000100",
                             4110 when "10111110000101",
                             4110 when "10111110000110",
                             4109 when "10111110000111",
                             4109 when "10111110001000",
                             4109 when "10111110001001",
                             4108 when "10111110001010",
                             4108 when "10111110001011",
                             4108 when "10111110001100",
                             4107 when "10111110001101",
                             4107 when "10111110001110",
                             4107 when "10111110001111",
                             4106 when "10111110010000",
                             4106 when "10111110010001",
                             4106 when "10111110010010",
                             4105 when "10111110010011",
                             4105 when "10111110010100",
                             4105 when "10111110010101",
                             4104 when "10111110010110",
                             4104 when "10111110010111",
                             4104 when "10111110011000",
                             4103 when "10111110011001",
                             4103 when "10111110011010",
                             4103 when "10111110011011",
                             4102 when "10111110011100",
                             4102 when "10111110011101",
                             4102 when "10111110011110",
                             4101 when "10111110011111",
                             4101 when "10111110100000",
                             4101 when "10111110100001",
                             4100 when "10111110100010",
                             4100 when "10111110100011",
                             4100 when "10111110100100",
                             4099 when "10111110100101",
                             4099 when "10111110100110",
                             4099 when "10111110100111",
                             4098 when "10111110101000",
                             4098 when "10111110101001",
                             4098 when "10111110101010",
                             4097 when "10111110101011",
                             4097 when "10111110101100",
                             4097 when "10111110101101",
                             4096 when "10111110101110",
                             4096 when "10111110101111",
                             4096 when "10111110110000",
                             4095 when "10111110110001",
                             4095 when "10111110110010",
                             4095 when "10111110110011",
                             4094 when "10111110110100",
                             4094 when "10111110110101",
                             4094 when "10111110110110",
                             4093 when "10111110110111",
                             4093 when "10111110111000",
                             4093 when "10111110111001",
                             4092 when "10111110111010",
                             4092 when "10111110111011",
                             4092 when "10111110111100",
                             4091 when "10111110111101",
                             4091 when "10111110111110",
                             4091 when "10111110111111",
                             4090 when "10111111000000",
                             4090 when "10111111000001",
                             4090 when "10111111000010",
                             4089 when "10111111000011",
                             4089 when "10111111000100",
                             4089 when "10111111000101",
                             4088 when "10111111000110",
                             4088 when "10111111000111",
                             4088 when "10111111001000",
                             4087 when "10111111001001",
                             4087 when "10111111001010",
                             4087 when "10111111001011",
                             4086 when "10111111001100",
                             4086 when "10111111001101",
                             4086 when "10111111001110",
                             4085 when "10111111001111",
                             4085 when "10111111010000",
                             4085 when "10111111010001",
                             4084 when "10111111010010",
                             4084 when "10111111010011",
                             4084 when "10111111010100",
                             4083 when "10111111010101",
                             4083 when "10111111010110",
                             4083 when "10111111010111",
                             4082 when "10111111011000",
                             4082 when "10111111011001",
                             4082 when "10111111011010",
                             4081 when "10111111011011",
                             4081 when "10111111011100",
                             4081 when "10111111011101",
                             4080 when "10111111011110",
                             4080 when "10111111011111",
                             4080 when "10111111100000",
                             4079 when "10111111100001",
                             4079 when "10111111100010",
                             4079 when "10111111100011",
                             4078 when "10111111100100",
                             4078 when "10111111100101",
                             4078 when "10111111100110",
                             4077 when "10111111100111",
                             4077 when "10111111101000",
                             4077 when "10111111101001",
                             4076 when "10111111101010",
                             4076 when "10111111101011",
                             4076 when "10111111101100",
                             4075 when "10111111101101",
                             4075 when "10111111101110",
                             4075 when "10111111101111",
                             4074 when "10111111110000",
                             4074 when "10111111110001",
                             4074 when "10111111110010",
                             4073 when "10111111110011",
                             4073 when "10111111110100",
                             4073 when "10111111110101",
                             4072 when "10111111110110",
                             4072 when "10111111110111",
                             4072 when "10111111111000",
                             4071 when "10111111111001",
                             4071 when "10111111111010",
                             4071 when "10111111111011",
                             4070 when "10111111111100",
                             4070 when "10111111111101",
                             4070 when "10111111111110",
                             4069 when "10111111111111",
                             4069 when "11000000000000",
                             4069 when "11000000000001",
                             4068 when "11000000000010",
                             4068 when "11000000000011",
                             4068 when "11000000000100",
                             4067 when "11000000000101",
                             4067 when "11000000000110",
                             4067 when "11000000000111",
                             4066 when "11000000001000",
                             4066 when "11000000001001",
                             4066 when "11000000001010",
                             4065 when "11000000001011",
                             4065 when "11000000001100",
                             4065 when "11000000001101",
                             4064 when "11000000001110",
                             4064 when "11000000001111",
                             4064 when "11000000010000",
                             4063 when "11000000010001",
                             4063 when "11000000010010",
                             4063 when "11000000010011",
                             4062 when "11000000010100",
                             4062 when "11000000010101",
                             4062 when "11000000010110",
                             4061 when "11000000010111",
                             4061 when "11000000011000",
                             4061 when "11000000011001",
                             4060 when "11000000011010",
                             4060 when "11000000011011",
                             4060 when "11000000011100",
                             4059 when "11000000011101",
                             4059 when "11000000011110",
                             4059 when "11000000011111",
                             4058 when "11000000100000",
                             4058 when "11000000100001",
                             4058 when "11000000100010",
                             4057 when "11000000100011",
                             4057 when "11000000100100",
                             4057 when "11000000100101",
                             4056 when "11000000100110",
                             4056 when "11000000100111",
                             4056 when "11000000101000",
                             4055 when "11000000101001",
                             4055 when "11000000101010",
                             4055 when "11000000101011",
                             4054 when "11000000101100",
                             4054 when "11000000101101",
                             4054 when "11000000101110",
                             4054 when "11000000101111",
                             4053 when "11000000110000",
                             4053 when "11000000110001",
                             4053 when "11000000110010",
                             4052 when "11000000110011",
                             4052 when "11000000110100",
                             4052 when "11000000110101",
                             4051 when "11000000110110",
                             4051 when "11000000110111",
                             4051 when "11000000111000",
                             4050 when "11000000111001",
                             4050 when "11000000111010",
                             4050 when "11000000111011",
                             4049 when "11000000111100",
                             4049 when "11000000111101",
                             4049 when "11000000111110",
                             4048 when "11000000111111",
                             4048 when "11000001000000",
                             4048 when "11000001000001",
                             4047 when "11000001000010",
                             4047 when "11000001000011",
                             4047 when "11000001000100",
                             4046 when "11000001000101",
                             4046 when "11000001000110",
                             4046 when "11000001000111",
                             4045 when "11000001001000",
                             4045 when "11000001001001",
                             4045 when "11000001001010",
                             4044 when "11000001001011",
                             4044 when "11000001001100",
                             4044 when "11000001001101",
                             4043 when "11000001001110",
                             4043 when "11000001001111",
                             4043 when "11000001010000",
                             4042 when "11000001010001",
                             4042 when "11000001010010",
                             4042 when "11000001010011",
                             4041 when "11000001010100",
                             4041 when "11000001010101",
                             4041 when "11000001010110",
                             4040 when "11000001010111",
                             4040 when "11000001011000",
                             4040 when "11000001011001",
                             4039 when "11000001011010",
                             4039 when "11000001011011",
                             4039 when "11000001011100",
                             4038 when "11000001011101",
                             4038 when "11000001011110",
                             4038 when "11000001011111",
                             4037 when "11000001100000",
                             4037 when "11000001100001",
                             4037 when "11000001100010",
                             4036 when "11000001100011",
                             4036 when "11000001100100",
                             4036 when "11000001100101",
                             4036 when "11000001100110",
                             4035 when "11000001100111",
                             4035 when "11000001101000",
                             4035 when "11000001101001",
                             4034 when "11000001101010",
                             4034 when "11000001101011",
                             4034 when "11000001101100",
                             4033 when "11000001101101",
                             4033 when "11000001101110",
                             4033 when "11000001101111",
                             4032 when "11000001110000",
                             4032 when "11000001110001",
                             4032 when "11000001110010",
                             4031 when "11000001110011",
                             4031 when "11000001110100",
                             4031 when "11000001110101",
                             4030 when "11000001110110",
                             4030 when "11000001110111",
                             4030 when "11000001111000",
                             4029 when "11000001111001",
                             4029 when "11000001111010",
                             4029 when "11000001111011",
                             4028 when "11000001111100",
                             4028 when "11000001111101",
                             4028 when "11000001111110",
                             4027 when "11000001111111",
                             4027 when "11000010000000",
                             4027 when "11000010000001",
                             4026 when "11000010000010",
                             4026 when "11000010000011",
                             4026 when "11000010000100",
                             4025 when "11000010000101",
                             4025 when "11000010000110",
                             4025 when "11000010000111",
                             4024 when "11000010001000",
                             4024 when "11000010001001",
                             4024 when "11000010001010",
                             4023 when "11000010001011",
                             4023 when "11000010001100",
                             4023 when "11000010001101",
                             4023 when "11000010001110",
                             4022 when "11000010001111",
                             4022 when "11000010010000",
                             4022 when "11000010010001",
                             4021 when "11000010010010",
                             4021 when "11000010010011",
                             4021 when "11000010010100",
                             4020 when "11000010010101",
                             4020 when "11000010010110",
                             4020 when "11000010010111",
                             4019 when "11000010011000",
                             4019 when "11000010011001",
                             4019 when "11000010011010",
                             4018 when "11000010011011",
                             4018 when "11000010011100",
                             4018 when "11000010011101",
                             4017 when "11000010011110",
                             4017 when "11000010011111",
                             4017 when "11000010100000",
                             4016 when "11000010100001",
                             4016 when "11000010100010",
                             4016 when "11000010100011",
                             4015 when "11000010100100",
                             4015 when "11000010100101",
                             4015 when "11000010100110",
                             4014 when "11000010100111",
                             4014 when "11000010101000",
                             4014 when "11000010101001",
                             4013 when "11000010101010",
                             4013 when "11000010101011",
                             4013 when "11000010101100",
                             4013 when "11000010101101",
                             4012 when "11000010101110",
                             4012 when "11000010101111",
                             4012 when "11000010110000",
                             4011 when "11000010110001",
                             4011 when "11000010110010",
                             4011 when "11000010110011",
                             4010 when "11000010110100",
                             4010 when "11000010110101",
                             4010 when "11000010110110",
                             4009 when "11000010110111",
                             4009 when "11000010111000",
                             4009 when "11000010111001",
                             4008 when "11000010111010",
                             4008 when "11000010111011",
                             4008 when "11000010111100",
                             4007 when "11000010111101",
                             4007 when "11000010111110",
                             4007 when "11000010111111",
                             4006 when "11000011000000",
                             4006 when "11000011000001",
                             4006 when "11000011000010",
                             4005 when "11000011000011",
                             4005 when "11000011000100",
                             4005 when "11000011000101",
                             4004 when "11000011000110",
                             4004 when "11000011000111",
                             4004 when "11000011001000",
                             4004 when "11000011001001",
                             4003 when "11000011001010",
                             4003 when "11000011001011",
                             4003 when "11000011001100",
                             4002 when "11000011001101",
                             4002 when "11000011001110",
                             4002 when "11000011001111",
                             4001 when "11000011010000",
                             4001 when "11000011010001",
                             4001 when "11000011010010",
                             4000 when "11000011010011",
                             4000 when "11000011010100",
                             4000 when "11000011010101",
                             3999 when "11000011010110",
                             3999 when "11000011010111",
                             3999 when "11000011011000",
                             3998 when "11000011011001",
                             3998 when "11000011011010",
                             3998 when "11000011011011",
                             3997 when "11000011011100",
                             3997 when "11000011011101",
                             3997 when "11000011011110",
                             3996 when "11000011011111",
                             3996 when "11000011100000",
                             3996 when "11000011100001",
                             3996 when "11000011100010",
                             3995 when "11000011100011",
                             3995 when "11000011100100",
                             3995 when "11000011100101",
                             3994 when "11000011100110",
                             3994 when "11000011100111",
                             3994 when "11000011101000",
                             3993 when "11000011101001",
                             3993 when "11000011101010",
                             3993 when "11000011101011",
                             3992 when "11000011101100",
                             3992 when "11000011101101",
                             3992 when "11000011101110",
                             3991 when "11000011101111",
                             3991 when "11000011110000",
                             3991 when "11000011110001",
                             3990 when "11000011110010",
                             3990 when "11000011110011",
                             3990 when "11000011110100",
                             3989 when "11000011110101",
                             3989 when "11000011110110",
                             3989 when "11000011110111",
                             3989 when "11000011111000",
                             3988 when "11000011111001",
                             3988 when "11000011111010",
                             3988 when "11000011111011",
                             3987 when "11000011111100",
                             3987 when "11000011111101",
                             3987 when "11000011111110",
                             3986 when "11000011111111",
                             3986 when "11000100000000",
                             3986 when "11000100000001",
                             3985 when "11000100000010",
                             3985 when "11000100000011",
                             3985 when "11000100000100",
                             3984 when "11000100000101",
                             3984 when "11000100000110",
                             3984 when "11000100000111",
                             3983 when "11000100001000",
                             3983 when "11000100001001",
                             3983 when "11000100001010",
                             3982 when "11000100001011",
                             3982 when "11000100001100",
                             3982 when "11000100001101",
                             3982 when "11000100001110",
                             3981 when "11000100001111",
                             3981 when "11000100010000",
                             3981 when "11000100010001",
                             3980 when "11000100010010",
                             3980 when "11000100010011",
                             3980 when "11000100010100",
                             3979 when "11000100010101",
                             3979 when "11000100010110",
                             3979 when "11000100010111",
                             3978 when "11000100011000",
                             3978 when "11000100011001",
                             3978 when "11000100011010",
                             3977 when "11000100011011",
                             3977 when "11000100011100",
                             3977 when "11000100011101",
                             3976 when "11000100011110",
                             3976 when "11000100011111",
                             3976 when "11000100100000",
                             3976 when "11000100100001",
                             3975 when "11000100100010",
                             3975 when "11000100100011",
                             3975 when "11000100100100",
                             3974 when "11000100100101",
                             3974 when "11000100100110",
                             3974 when "11000100100111",
                             3973 when "11000100101000",
                             3973 when "11000100101001",
                             3973 when "11000100101010",
                             3972 when "11000100101011",
                             3972 when "11000100101100",
                             3972 when "11000100101101",
                             3971 when "11000100101110",
                             3971 when "11000100101111",
                             3971 when "11000100110000",
                             3970 when "11000100110001",
                             3970 when "11000100110010",
                             3970 when "11000100110011",
                             3970 when "11000100110100",
                             3969 when "11000100110101",
                             3969 when "11000100110110",
                             3969 when "11000100110111",
                             3968 when "11000100111000",
                             3968 when "11000100111001",
                             3968 when "11000100111010",
                             3967 when "11000100111011",
                             3967 when "11000100111100",
                             3967 when "11000100111101",
                             3966 when "11000100111110",
                             3966 when "11000100111111",
                             3966 when "11000101000000",
                             3965 when "11000101000001",
                             3965 when "11000101000010",
                             3965 when "11000101000011",
                             3964 when "11000101000100",
                             3964 when "11000101000101",
                             3964 when "11000101000110",
                             3964 when "11000101000111",
                             3963 when "11000101001000",
                             3963 when "11000101001001",
                             3963 when "11000101001010",
                             3962 when "11000101001011",
                             3962 when "11000101001100",
                             3962 when "11000101001101",
                             3961 when "11000101001110",
                             3961 when "11000101001111",
                             3961 when "11000101010000",
                             3960 when "11000101010001",
                             3960 when "11000101010010",
                             3960 when "11000101010011",
                             3959 when "11000101010100",
                             3959 when "11000101010101",
                             3959 when "11000101010110",
                             3959 when "11000101010111",
                             3958 when "11000101011000",
                             3958 when "11000101011001",
                             3958 when "11000101011010",
                             3957 when "11000101011011",
                             3957 when "11000101011100",
                             3957 when "11000101011101",
                             3956 when "11000101011110",
                             3956 when "11000101011111",
                             3956 when "11000101100000",
                             3955 when "11000101100001",
                             3955 when "11000101100010",
                             3955 when "11000101100011",
                             3954 when "11000101100100",
                             3954 when "11000101100101",
                             3954 when "11000101100110",
                             3954 when "11000101100111",
                             3953 when "11000101101000",
                             3953 when "11000101101001",
                             3953 when "11000101101010",
                             3952 when "11000101101011",
                             3952 when "11000101101100",
                             3952 when "11000101101101",
                             3951 when "11000101101110",
                             3951 when "11000101101111",
                             3951 when "11000101110000",
                             3950 when "11000101110001",
                             3950 when "11000101110010",
                             3950 when "11000101110011",
                             3949 when "11000101110100",
                             3949 when "11000101110101",
                             3949 when "11000101110110",
                             3949 when "11000101110111",
                             3948 when "11000101111000",
                             3948 when "11000101111001",
                             3948 when "11000101111010",
                             3947 when "11000101111011",
                             3947 when "11000101111100",
                             3947 when "11000101111101",
                             3946 when "11000101111110",
                             3946 when "11000101111111",
                             3946 when "11000110000000",
                             3945 when "11000110000001",
                             3945 when "11000110000010",
                             3945 when "11000110000011",
                             3944 when "11000110000100",
                             3944 when "11000110000101",
                             3944 when "11000110000110",
                             3944 when "11000110000111",
                             3943 when "11000110001000",
                             3943 when "11000110001001",
                             3943 when "11000110001010",
                             3942 when "11000110001011",
                             3942 when "11000110001100",
                             3942 when "11000110001101",
                             3941 when "11000110001110",
                             3941 when "11000110001111",
                             3941 when "11000110010000",
                             3940 when "11000110010001",
                             3940 when "11000110010010",
                             3940 when "11000110010011",
                             3939 when "11000110010100",
                             3939 when "11000110010101",
                             3939 when "11000110010110",
                             3939 when "11000110010111",
                             3938 when "11000110011000",
                             3938 when "11000110011001",
                             3938 when "11000110011010",
                             3937 when "11000110011011",
                             3937 when "11000110011100",
                             3937 when "11000110011101",
                             3936 when "11000110011110",
                             3936 when "11000110011111",
                             3936 when "11000110100000",
                             3935 when "11000110100001",
                             3935 when "11000110100010",
                             3935 when "11000110100011",
                             3935 when "11000110100100",
                             3934 when "11000110100101",
                             3934 when "11000110100110",
                             3934 when "11000110100111",
                             3933 when "11000110101000",
                             3933 when "11000110101001",
                             3933 when "11000110101010",
                             3932 when "11000110101011",
                             3932 when "11000110101100",
                             3932 when "11000110101101",
                             3931 when "11000110101110",
                             3931 when "11000110101111",
                             3931 when "11000110110000",
                             3931 when "11000110110001",
                             3930 when "11000110110010",
                             3930 when "11000110110011",
                             3930 when "11000110110100",
                             3929 when "11000110110101",
                             3929 when "11000110110110",
                             3929 when "11000110110111",
                             3928 when "11000110111000",
                             3928 when "11000110111001",
                             3928 when "11000110111010",
                             3927 when "11000110111011",
                             3927 when "11000110111100",
                             3927 when "11000110111101",
                             3926 when "11000110111110",
                             3926 when "11000110111111",
                             3926 when "11000111000000",
                             3926 when "11000111000001",
                             3925 when "11000111000010",
                             3925 when "11000111000011",
                             3925 when "11000111000100",
                             3924 when "11000111000101",
                             3924 when "11000111000110",
                             3924 when "11000111000111",
                             3923 when "11000111001000",
                             3923 when "11000111001001",
                             3923 when "11000111001010",
                             3922 when "11000111001011",
                             3922 when "11000111001100",
                             3922 when "11000111001101",
                             3922 when "11000111001110",
                             3921 when "11000111001111",
                             3921 when "11000111010000",
                             3921 when "11000111010001",
                             3920 when "11000111010010",
                             3920 when "11000111010011",
                             3920 when "11000111010100",
                             3919 when "11000111010101",
                             3919 when "11000111010110",
                             3919 when "11000111010111",
                             3918 when "11000111011000",
                             3918 when "11000111011001",
                             3918 when "11000111011010",
                             3918 when "11000111011011",
                             3917 when "11000111011100",
                             3917 when "11000111011101",
                             3917 when "11000111011110",
                             3916 when "11000111011111",
                             3916 when "11000111100000",
                             3916 when "11000111100001",
                             3915 when "11000111100010",
                             3915 when "11000111100011",
                             3915 when "11000111100100",
                             3915 when "11000111100101",
                             3914 when "11000111100110",
                             3914 when "11000111100111",
                             3914 when "11000111101000",
                             3913 when "11000111101001",
                             3913 when "11000111101010",
                             3913 when "11000111101011",
                             3912 when "11000111101100",
                             3912 when "11000111101101",
                             3912 when "11000111101110",
                             3911 when "11000111101111",
                             3911 when "11000111110000",
                             3911 when "11000111110001",
                             3911 when "11000111110010",
                             3910 when "11000111110011",
                             3910 when "11000111110100",
                             3910 when "11000111110101",
                             3909 when "11000111110110",
                             3909 when "11000111110111",
                             3909 when "11000111111000",
                             3908 when "11000111111001",
                             3908 when "11000111111010",
                             3908 when "11000111111011",
                             3907 when "11000111111100",
                             3907 when "11000111111101",
                             3907 when "11000111111110",
                             3907 when "11000111111111",
                             3906 when "11001000000000",
                             3906 when "11001000000001",
                             3906 when "11001000000010",
                             3905 when "11001000000011",
                             3905 when "11001000000100",
                             3905 when "11001000000101",
                             3904 when "11001000000110",
                             3904 when "11001000000111",
                             3904 when "11001000001000",
                             3904 when "11001000001001",
                             3903 when "11001000001010",
                             3903 when "11001000001011",
                             3903 when "11001000001100",
                             3902 when "11001000001101",
                             3902 when "11001000001110",
                             3902 when "11001000001111",
                             3901 when "11001000010000",
                             3901 when "11001000010001",
                             3901 when "11001000010010",
                             3900 when "11001000010011",
                             3900 when "11001000010100",
                             3900 when "11001000010101",
                             3900 when "11001000010110",
                             3899 when "11001000010111",
                             3899 when "11001000011000",
                             3899 when "11001000011001",
                             3898 when "11001000011010",
                             3898 when "11001000011011",
                             3898 when "11001000011100",
                             3897 when "11001000011101",
                             3897 when "11001000011110",
                             3897 when "11001000011111",
                             3897 when "11001000100000",
                             3896 when "11001000100001",
                             3896 when "11001000100010",
                             3896 when "11001000100011",
                             3895 when "11001000100100",
                             3895 when "11001000100101",
                             3895 when "11001000100110",
                             3894 when "11001000100111",
                             3894 when "11001000101000",
                             3894 when "11001000101001",
                             3893 when "11001000101010",
                             3893 when "11001000101011",
                             3893 when "11001000101100",
                             3893 when "11001000101101",
                             3892 when "11001000101110",
                             3892 when "11001000101111",
                             3892 when "11001000110000",
                             3891 when "11001000110001",
                             3891 when "11001000110010",
                             3891 when "11001000110011",
                             3890 when "11001000110100",
                             3890 when "11001000110101",
                             3890 when "11001000110110",
                             3890 when "11001000110111",
                             3889 when "11001000111000",
                             3889 when "11001000111001",
                             3889 when "11001000111010",
                             3888 when "11001000111011",
                             3888 when "11001000111100",
                             3888 when "11001000111101",
                             3887 when "11001000111110",
                             3887 when "11001000111111",
                             3887 when "11001001000000",
                             3887 when "11001001000001",
                             3886 when "11001001000010",
                             3886 when "11001001000011",
                             3886 when "11001001000100",
                             3885 when "11001001000101",
                             3885 when "11001001000110",
                             3885 when "11001001000111",
                             3884 when "11001001001000",
                             3884 when "11001001001001",
                             3884 when "11001001001010",
                             3883 when "11001001001011",
                             3883 when "11001001001100",
                             3883 when "11001001001101",
                             3883 when "11001001001110",
                             3882 when "11001001001111",
                             3882 when "11001001010000",
                             3882 when "11001001010001",
                             3881 when "11001001010010",
                             3881 when "11001001010011",
                             3881 when "11001001010100",
                             3880 when "11001001010101",
                             3880 when "11001001010110",
                             3880 when "11001001010111",
                             3880 when "11001001011000",
                             3879 when "11001001011001",
                             3879 when "11001001011010",
                             3879 when "11001001011011",
                             3878 when "11001001011100",
                             3878 when "11001001011101",
                             3878 when "11001001011110",
                             3877 when "11001001011111",
                             3877 when "11001001100000",
                             3877 when "11001001100001",
                             3877 when "11001001100010",
                             3876 when "11001001100011",
                             3876 when "11001001100100",
                             3876 when "11001001100101",
                             3875 when "11001001100110",
                             3875 when "11001001100111",
                             3875 when "11001001101000",
                             3874 when "11001001101001",
                             3874 when "11001001101010",
                             3874 when "11001001101011",
                             3874 when "11001001101100",
                             3873 when "11001001101101",
                             3873 when "11001001101110",
                             3873 when "11001001101111",
                             3872 when "11001001110000",
                             3872 when "11001001110001",
                             3872 when "11001001110010",
                             3871 when "11001001110011",
                             3871 when "11001001110100",
                             3871 when "11001001110101",
                             3871 when "11001001110110",
                             3870 when "11001001110111",
                             3870 when "11001001111000",
                             3870 when "11001001111001",
                             3869 when "11001001111010",
                             3869 when "11001001111011",
                             3869 when "11001001111100",
                             3868 when "11001001111101",
                             3868 when "11001001111110",
                             3868 when "11001001111111",
                             3868 when "11001010000000",
                             3867 when "11001010000001",
                             3867 when "11001010000010",
                             3867 when "11001010000011",
                             3866 when "11001010000100",
                             3866 when "11001010000101",
                             3866 when "11001010000110",
                             3865 when "11001010000111",
                             3865 when "11001010001000",
                             3865 when "11001010001001",
                             3865 when "11001010001010",
                             3864 when "11001010001011",
                             3864 when "11001010001100",
                             3864 when "11001010001101",
                             3863 when "11001010001110",
                             3863 when "11001010001111",
                             3863 when "11001010010000",
                             3862 when "11001010010001",
                             3862 when "11001010010010",
                             3862 when "11001010010011",
                             3862 when "11001010010100",
                             3861 when "11001010010101",
                             3861 when "11001010010110",
                             3861 when "11001010010111",
                             3860 when "11001010011000",
                             3860 when "11001010011001",
                             3860 when "11001010011010",
                             3860 when "11001010011011",
                             3859 when "11001010011100",
                             3859 when "11001010011101",
                             3859 when "11001010011110",
                             3858 when "11001010011111",
                             3858 when "11001010100000",
                             3858 when "11001010100001",
                             3857 when "11001010100010",
                             3857 when "11001010100011",
                             3857 when "11001010100100",
                             3857 when "11001010100101",
                             3856 when "11001010100110",
                             3856 when "11001010100111",
                             3856 when "11001010101000",
                             3855 when "11001010101001",
                             3855 when "11001010101010",
                             3855 when "11001010101011",
                             3854 when "11001010101100",
                             3854 when "11001010101101",
                             3854 when "11001010101110",
                             3854 when "11001010101111",
                             3853 when "11001010110000",
                             3853 when "11001010110001",
                             3853 when "11001010110010",
                             3852 when "11001010110011",
                             3852 when "11001010110100",
                             3852 when "11001010110101",
                             3851 when "11001010110110",
                             3851 when "11001010110111",
                             3851 when "11001010111000",
                             3851 when "11001010111001",
                             3850 when "11001010111010",
                             3850 when "11001010111011",
                             3850 when "11001010111100",
                             3849 when "11001010111101",
                             3849 when "11001010111110",
                             3849 when "11001010111111",
                             3849 when "11001011000000",
                             3848 when "11001011000001",
                             3848 when "11001011000010",
                             3848 when "11001011000011",
                             3847 when "11001011000100",
                             3847 when "11001011000101",
                             3847 when "11001011000110",
                             3846 when "11001011000111",
                             3846 when "11001011001000",
                             3846 when "11001011001001",
                             3846 when "11001011001010",
                             3845 when "11001011001011",
                             3845 when "11001011001100",
                             3845 when "11001011001101",
                             3844 when "11001011001110",
                             3844 when "11001011001111",
                             3844 when "11001011010000",
                             3843 when "11001011010001",
                             3843 when "11001011010010",
                             3843 when "11001011010011",
                             3843 when "11001011010100",
                             3842 when "11001011010101",
                             3842 when "11001011010110",
                             3842 when "11001011010111",
                             3841 when "11001011011000",
                             3841 when "11001011011001",
                             3841 when "11001011011010",
                             3841 when "11001011011011",
                             3840 when "11001011011100",
                             3840 when "11001011011101",
                             3840 when "11001011011110",
                             3839 when "11001011011111",
                             3839 when "11001011100000",
                             3839 when "11001011100001",
                             3838 when "11001011100010",
                             3838 when "11001011100011",
                             3838 when "11001011100100",
                             3838 when "11001011100101",
                             3837 when "11001011100110",
                             3837 when "11001011100111",
                             3837 when "11001011101000",
                             3836 when "11001011101001",
                             3836 when "11001011101010",
                             3836 when "11001011101011",
                             3836 when "11001011101100",
                             3835 when "11001011101101",
                             3835 when "11001011101110",
                             3835 when "11001011101111",
                             3834 when "11001011110000",
                             3834 when "11001011110001",
                             3834 when "11001011110010",
                             3833 when "11001011110011",
                             3833 when "11001011110100",
                             3833 when "11001011110101",
                             3833 when "11001011110110",
                             3832 when "11001011110111",
                             3832 when "11001011111000",
                             3832 when "11001011111001",
                             3831 when "11001011111010",
                             3831 when "11001011111011",
                             3831 when "11001011111100",
                             3831 when "11001011111101",
                             3830 when "11001011111110",
                             3830 when "11001011111111",
                             3830 when "11001100000000",
                             3829 when "11001100000001",
                             3829 when "11001100000010",
                             3829 when "11001100000011",
                             3828 when "11001100000100",
                             3828 when "11001100000101",
                             3828 when "11001100000110",
                             3828 when "11001100000111",
                             3827 when "11001100001000",
                             3827 when "11001100001001",
                             3827 when "11001100001010",
                             3826 when "11001100001011",
                             3826 when "11001100001100",
                             3826 when "11001100001101",
                             3826 when "11001100001110",
                             3825 when "11001100001111",
                             3825 when "11001100010000",
                             3825 when "11001100010001",
                             3824 when "11001100010010",
                             3824 when "11001100010011",
                             3824 when "11001100010100",
                             3824 when "11001100010101",
                             3823 when "11001100010110",
                             3823 when "11001100010111",
                             3823 when "11001100011000",
                             3822 when "11001100011001",
                             3822 when "11001100011010",
                             3822 when "11001100011011",
                             3821 when "11001100011100",
                             3821 when "11001100011101",
                             3821 when "11001100011110",
                             3821 when "11001100011111",
                             3820 when "11001100100000",
                             3820 when "11001100100001",
                             3820 when "11001100100010",
                             3819 when "11001100100011",
                             3819 when "11001100100100",
                             3819 when "11001100100101",
                             3819 when "11001100100110",
                             3818 when "11001100100111",
                             3818 when "11001100101000",
                             3818 when "11001100101001",
                             3817 when "11001100101010",
                             3817 when "11001100101011",
                             3817 when "11001100101100",
                             3817 when "11001100101101",
                             3816 when "11001100101110",
                             3816 when "11001100101111",
                             3816 when "11001100110000",
                             3815 when "11001100110001",
                             3815 when "11001100110010",
                             3815 when "11001100110011",
                             3814 when "11001100110100",
                             3814 when "11001100110101",
                             3814 when "11001100110110",
                             3814 when "11001100110111",
                             3813 when "11001100111000",
                             3813 when "11001100111001",
                             3813 when "11001100111010",
                             3812 when "11001100111011",
                             3812 when "11001100111100",
                             3812 when "11001100111101",
                             3812 when "11001100111110",
                             3811 when "11001100111111",
                             3811 when "11001101000000",
                             3811 when "11001101000001",
                             3810 when "11001101000010",
                             3810 when "11001101000011",
                             3810 when "11001101000100",
                             3810 when "11001101000101",
                             3809 when "11001101000110",
                             3809 when "11001101000111",
                             3809 when "11001101001000",
                             3808 when "11001101001001",
                             3808 when "11001101001010",
                             3808 when "11001101001011",
                             3807 when "11001101001100",
                             3807 when "11001101001101",
                             3807 when "11001101001110",
                             3807 when "11001101001111",
                             3806 when "11001101010000",
                             3806 when "11001101010001",
                             3806 when "11001101010010",
                             3805 when "11001101010011",
                             3805 when "11001101010100",
                             3805 when "11001101010101",
                             3805 when "11001101010110",
                             3804 when "11001101010111",
                             3804 when "11001101011000",
                             3804 when "11001101011001",
                             3803 when "11001101011010",
                             3803 when "11001101011011",
                             3803 when "11001101011100",
                             3803 when "11001101011101",
                             3802 when "11001101011110",
                             3802 when "11001101011111",
                             3802 when "11001101100000",
                             3801 when "11001101100001",
                             3801 when "11001101100010",
                             3801 when "11001101100011",
                             3801 when "11001101100100",
                             3800 when "11001101100101",
                             3800 when "11001101100110",
                             3800 when "11001101100111",
                             3799 when "11001101101000",
                             3799 when "11001101101001",
                             3799 when "11001101101010",
                             3799 when "11001101101011",
                             3798 when "11001101101100",
                             3798 when "11001101101101",
                             3798 when "11001101101110",
                             3797 when "11001101101111",
                             3797 when "11001101110000",
                             3797 when "11001101110001",
                             3797 when "11001101110010",
                             3796 when "11001101110011",
                             3796 when "11001101110100",
                             3796 when "11001101110101",
                             3795 when "11001101110110",
                             3795 when "11001101110111",
                             3795 when "11001101111000",
                             3794 when "11001101111001",
                             3794 when "11001101111010",
                             3794 when "11001101111011",
                             3794 when "11001101111100",
                             3793 when "11001101111101",
                             3793 when "11001101111110",
                             3793 when "11001101111111",
                             3792 when "11001110000000",
                             3792 when "11001110000001",
                             3792 when "11001110000010",
                             3792 when "11001110000011",
                             3791 when "11001110000100",
                             3791 when "11001110000101",
                             3791 when "11001110000110",
                             3790 when "11001110000111",
                             3790 when "11001110001000",
                             3790 when "11001110001001",
                             3790 when "11001110001010",
                             3789 when "11001110001011",
                             3789 when "11001110001100",
                             3789 when "11001110001101",
                             3788 when "11001110001110",
                             3788 when "11001110001111",
                             3788 when "11001110010000",
                             3788 when "11001110010001",
                             3787 when "11001110010010",
                             3787 when "11001110010011",
                             3787 when "11001110010100",
                             3786 when "11001110010101",
                             3786 when "11001110010110",
                             3786 when "11001110010111",
                             3786 when "11001110011000",
                             3785 when "11001110011001",
                             3785 when "11001110011010",
                             3785 when "11001110011011",
                             3784 when "11001110011100",
                             3784 when "11001110011101",
                             3784 when "11001110011110",
                             3784 when "11001110011111",
                             3783 when "11001110100000",
                             3783 when "11001110100001",
                             3783 when "11001110100010",
                             3782 when "11001110100011",
                             3782 when "11001110100100",
                             3782 when "11001110100101",
                             3782 when "11001110100110",
                             3781 when "11001110100111",
                             3781 when "11001110101000",
                             3781 when "11001110101001",
                             3780 when "11001110101010",
                             3780 when "11001110101011",
                             3780 when "11001110101100",
                             3780 when "11001110101101",
                             3779 when "11001110101110",
                             3779 when "11001110101111",
                             3779 when "11001110110000",
                             3778 when "11001110110001",
                             3778 when "11001110110010",
                             3778 when "11001110110011",
                             3778 when "11001110110100",
                             3777 when "11001110110101",
                             3777 when "11001110110110",
                             3777 when "11001110110111",
                             3776 when "11001110111000",
                             3776 when "11001110111001",
                             3776 when "11001110111010",
                             3776 when "11001110111011",
                             3775 when "11001110111100",
                             3775 when "11001110111101",
                             3775 when "11001110111110",
                             3774 when "11001110111111",
                             3774 when "11001111000000",
                             3774 when "11001111000001",
                             3774 when "11001111000010",
                             3773 when "11001111000011",
                             3773 when "11001111000100",
                             3773 when "11001111000101",
                             3772 when "11001111000110",
                             3772 when "11001111000111",
                             3772 when "11001111001000",
                             3772 when "11001111001001",
                             3771 when "11001111001010",
                             3771 when "11001111001011",
                             3771 when "11001111001100",
                             3770 when "11001111001101",
                             3770 when "11001111001110",
                             3770 when "11001111001111",
                             3770 when "11001111010000",
                             3769 when "11001111010001",
                             3769 when "11001111010010",
                             3769 when "11001111010011",
                             3768 when "11001111010100",
                             3768 when "11001111010101",
                             3768 when "11001111010110",
                             3768 when "11001111010111",
                             3767 when "11001111011000",
                             3767 when "11001111011001",
                             3767 when "11001111011010",
                             3766 when "11001111011011",
                             3766 when "11001111011100",
                             3766 when "11001111011101",
                             3766 when "11001111011110",
                             3765 when "11001111011111",
                             3765 when "11001111100000",
                             3765 when "11001111100001",
                             3764 when "11001111100010",
                             3764 when "11001111100011",
                             3764 when "11001111100100",
                             3764 when "11001111100101",
                             3763 when "11001111100110",
                             3763 when "11001111100111",
                             3763 when "11001111101000",
                             3763 when "11001111101001",
                             3762 when "11001111101010",
                             3762 when "11001111101011",
                             3762 when "11001111101100",
                             3761 when "11001111101101",
                             3761 when "11001111101110",
                             3761 when "11001111101111",
                             3761 when "11001111110000",
                             3760 when "11001111110001",
                             3760 when "11001111110010",
                             3760 when "11001111110011",
                             3759 when "11001111110100",
                             3759 when "11001111110101",
                             3759 when "11001111110110",
                             3759 when "11001111110111",
                             3758 when "11001111111000",
                             3758 when "11001111111001",
                             3758 when "11001111111010",
                             3757 when "11001111111011",
                             3757 when "11001111111100",
                             3757 when "11001111111101",
                             3757 when "11001111111110",
                             3756 when "11001111111111",
                             3756 when "11010000000000",
                             3756 when "11010000000001",
                             3755 when "11010000000010",
                             3755 when "11010000000011",
                             3755 when "11010000000100",
                             3755 when "11010000000101",
                             3754 when "11010000000110",
                             3754 when "11010000000111",
                             3754 when "11010000001000",
                             3753 when "11010000001001",
                             3753 when "11010000001010",
                             3753 when "11010000001011",
                             3753 when "11010000001100",
                             3752 when "11010000001101",
                             3752 when "11010000001110",
                             3752 when "11010000001111",
                             3752 when "11010000010000",
                             3751 when "11010000010001",
                             3751 when "11010000010010",
                             3751 when "11010000010011",
                             3750 when "11010000010100",
                             3750 when "11010000010101",
                             3750 when "11010000010110",
                             3750 when "11010000010111",
                             3749 when "11010000011000",
                             3749 when "11010000011001",
                             3749 when "11010000011010",
                             3748 when "11010000011011",
                             3748 when "11010000011100",
                             3748 when "11010000011101",
                             3748 when "11010000011110",
                             3747 when "11010000011111",
                             3747 when "11010000100000",
                             3747 when "11010000100001",
                             3746 when "11010000100010",
                             3746 when "11010000100011",
                             3746 when "11010000100100",
                             3746 when "11010000100101",
                             3745 when "11010000100110",
                             3745 when "11010000100111",
                             3745 when "11010000101000",
                             3744 when "11010000101001",
                             3744 when "11010000101010",
                             3744 when "11010000101011",
                             3744 when "11010000101100",
                             3743 when "11010000101101",
                             3743 when "11010000101110",
                             3743 when "11010000101111",
                             3743 when "11010000110000",
                             3742 when "11010000110001",
                             3742 when "11010000110010",
                             3742 when "11010000110011",
                             3741 when "11010000110100",
                             3741 when "11010000110101",
                             3741 when "11010000110110",
                             3741 when "11010000110111",
                             3740 when "11010000111000",
                             3740 when "11010000111001",
                             3740 when "11010000111010",
                             3739 when "11010000111011",
                             3739 when "11010000111100",
                             3739 when "11010000111101",
                             3739 when "11010000111110",
                             3738 when "11010000111111",
                             3738 when "11010001000000",
                             3738 when "11010001000001",
                             3737 when "11010001000010",
                             3737 when "11010001000011",
                             3737 when "11010001000100",
                             3737 when "11010001000101",
                             3736 when "11010001000110",
                             3736 when "11010001000111",
                             3736 when "11010001001000",
                             3736 when "11010001001001",
                             3735 when "11010001001010",
                             3735 when "11010001001011",
                             3735 when "11010001001100",
                             3734 when "11010001001101",
                             3734 when "11010001001110",
                             3734 when "11010001001111",
                             3734 when "11010001010000",
                             3733 when "11010001010001",
                             3733 when "11010001010010",
                             3733 when "11010001010011",
                             3732 when "11010001010100",
                             3732 when "11010001010101",
                             3732 when "11010001010110",
                             3732 when "11010001010111",
                             3731 when "11010001011000",
                             3731 when "11010001011001",
                             3731 when "11010001011010",
                             3731 when "11010001011011",
                             3730 when "11010001011100",
                             3730 when "11010001011101",
                             3730 when "11010001011110",
                             3729 when "11010001011111",
                             3729 when "11010001100000",
                             3729 when "11010001100001",
                             3729 when "11010001100010",
                             3728 when "11010001100011",
                             3728 when "11010001100100",
                             3728 when "11010001100101",
                             3727 when "11010001100110",
                             3727 when "11010001100111",
                             3727 when "11010001101000",
                             3727 when "11010001101001",
                             3726 when "11010001101010",
                             3726 when "11010001101011",
                             3726 when "11010001101100",
                             3726 when "11010001101101",
                             3725 when "11010001101110",
                             3725 when "11010001101111",
                             3725 when "11010001110000",
                             3724 when "11010001110001",
                             3724 when "11010001110010",
                             3724 when "11010001110011",
                             3724 when "11010001110100",
                             3723 when "11010001110101",
                             3723 when "11010001110110",
                             3723 when "11010001110111",
                             3722 when "11010001111000",
                             3722 when "11010001111001",
                             3722 when "11010001111010",
                             3722 when "11010001111011",
                             3721 when "11010001111100",
                             3721 when "11010001111101",
                             3721 when "11010001111110",
                             3721 when "11010001111111",
                             3720 when "11010010000000",
                             3720 when "11010010000001",
                             3720 when "11010010000010",
                             3719 when "11010010000011",
                             3719 when "11010010000100",
                             3719 when "11010010000101",
                             3719 when "11010010000110",
                             3718 when "11010010000111",
                             3718 when "11010010001000",
                             3718 when "11010010001001",
                             3717 when "11010010001010",
                             3717 when "11010010001011",
                             3717 when "11010010001100",
                             3717 when "11010010001101",
                             3716 when "11010010001110",
                             3716 when "11010010001111",
                             3716 when "11010010010000",
                             3716 when "11010010010001",
                             3715 when "11010010010010",
                             3715 when "11010010010011",
                             3715 when "11010010010100",
                             3714 when "11010010010101",
                             3714 when "11010010010110",
                             3714 when "11010010010111",
                             3714 when "11010010011000",
                             3713 when "11010010011001",
                             3713 when "11010010011010",
                             3713 when "11010010011011",
                             3713 when "11010010011100",
                             3712 when "11010010011101",
                             3712 when "11010010011110",
                             3712 when "11010010011111",
                             3711 when "11010010100000",
                             3711 when "11010010100001",
                             3711 when "11010010100010",
                             3711 when "11010010100011",
                             3710 when "11010010100100",
                             3710 when "11010010100101",
                             3710 when "11010010100110",
                             3709 when "11010010100111",
                             3709 when "11010010101000",
                             3709 when "11010010101001",
                             3709 when "11010010101010",
                             3708 when "11010010101011",
                             3708 when "11010010101100",
                             3708 when "11010010101101",
                             3708 when "11010010101110",
                             3707 when "11010010101111",
                             3707 when "11010010110000",
                             3707 when "11010010110001",
                             3706 when "11010010110010",
                             3706 when "11010010110011",
                             3706 when "11010010110100",
                             3706 when "11010010110101",
                             3705 when "11010010110110",
                             3705 when "11010010110111",
                             3705 when "11010010111000",
                             3705 when "11010010111001",
                             3704 when "11010010111010",
                             3704 when "11010010111011",
                             3704 when "11010010111100",
                             3703 when "11010010111101",
                             3703 when "11010010111110",
                             3703 when "11010010111111",
                             3703 when "11010011000000",
                             3702 when "11010011000001",
                             3702 when "11010011000010",
                             3702 when "11010011000011",
                             3702 when "11010011000100",
                             3701 when "11010011000101",
                             3701 when "11010011000110",
                             3701 when "11010011000111",
                             3700 when "11010011001000",
                             3700 when "11010011001001",
                             3700 when "11010011001010",
                             3700 when "11010011001011",
                             3699 when "11010011001100",
                             3699 when "11010011001101",
                             3699 when "11010011001110",
                             3698 when "11010011001111",
                             3698 when "11010011010000",
                             3698 when "11010011010001",
                             3698 when "11010011010010",
                             3697 when "11010011010011",
                             3697 when "11010011010100",
                             3697 when "11010011010101",
                             3697 when "11010011010110",
                             3696 when "11010011010111",
                             3696 when "11010011011000",
                             3696 when "11010011011001",
                             3695 when "11010011011010",
                             3695 when "11010011011011",
                             3695 when "11010011011100",
                             3695 when "11010011011101",
                             3694 when "11010011011110",
                             3694 when "11010011011111",
                             3694 when "11010011100000",
                             3694 when "11010011100001",
                             3693 when "11010011100010",
                             3693 when "11010011100011",
                             3693 when "11010011100100",
                             3692 when "11010011100101",
                             3692 when "11010011100110",
                             3692 when "11010011100111",
                             3692 when "11010011101000",
                             3691 when "11010011101001",
                             3691 when "11010011101010",
                             3691 when "11010011101011",
                             3691 when "11010011101100",
                             3690 when "11010011101101",
                             3690 when "11010011101110",
                             3690 when "11010011101111",
                             3689 when "11010011110000",
                             3689 when "11010011110001",
                             3689 when "11010011110010",
                             3689 when "11010011110011",
                             3688 when "11010011110100",
                             3688 when "11010011110101",
                             3688 when "11010011110110",
                             3688 when "11010011110111",
                             3687 when "11010011111000",
                             3687 when "11010011111001",
                             3687 when "11010011111010",
                             3687 when "11010011111011",
                             3686 when "11010011111100",
                             3686 when "11010011111101",
                             3686 when "11010011111110",
                             3685 when "11010011111111",
                             3685 when "11010100000000",
                             3685 when "11010100000001",
                             3685 when "11010100000010",
                             3684 when "11010100000011",
                             3684 when "11010100000100",
                             3684 when "11010100000101",
                             3684 when "11010100000110",
                             3683 when "11010100000111",
                             3683 when "11010100001000",
                             3683 when "11010100001001",
                             3682 when "11010100001010",
                             3682 when "11010100001011",
                             3682 when "11010100001100",
                             3682 when "11010100001101",
                             3681 when "11010100001110",
                             3681 when "11010100001111",
                             3681 when "11010100010000",
                             3681 when "11010100010001",
                             3680 when "11010100010010",
                             3680 when "11010100010011",
                             3680 when "11010100010100",
                             3679 when "11010100010101",
                             3679 when "11010100010110",
                             3679 when "11010100010111",
                             3679 when "11010100011000",
                             3678 when "11010100011001",
                             3678 when "11010100011010",
                             3678 when "11010100011011",
                             3678 when "11010100011100",
                             3677 when "11010100011101",
                             3677 when "11010100011110",
                             3677 when "11010100011111",
                             3676 when "11010100100000",
                             3676 when "11010100100001",
                             3676 when "11010100100010",
                             3676 when "11010100100011",
                             3675 when "11010100100100",
                             3675 when "11010100100101",
                             3675 when "11010100100110",
                             3675 when "11010100100111",
                             3674 when "11010100101000",
                             3674 when "11010100101001",
                             3674 when "11010100101010",
                             3673 when "11010100101011",
                             3673 when "11010100101100",
                             3673 when "11010100101101",
                             3673 when "11010100101110",
                             3672 when "11010100101111",
                             3672 when "11010100110000",
                             3672 when "11010100110001",
                             3672 when "11010100110010",
                             3671 when "11010100110011",
                             3671 when "11010100110100",
                             3671 when "11010100110101",
                             3671 when "11010100110110",
                             3670 when "11010100110111",
                             3670 when "11010100111000",
                             3670 when "11010100111001",
                             3669 when "11010100111010",
                             3669 when "11010100111011",
                             3669 when "11010100111100",
                             3669 when "11010100111101",
                             3668 when "11010100111110",
                             3668 when "11010100111111",
                             3668 when "11010101000000",
                             3668 when "11010101000001",
                             3667 when "11010101000010",
                             3667 when "11010101000011",
                             3667 when "11010101000100",
                             3666 when "11010101000101",
                             3666 when "11010101000110",
                             3666 when "11010101000111",
                             3666 when "11010101001000",
                             3665 when "11010101001001",
                             3665 when "11010101001010",
                             3665 when "11010101001011",
                             3665 when "11010101001100",
                             3664 when "11010101001101",
                             3664 when "11010101001110",
                             3664 when "11010101001111",
                             3664 when "11010101010000",
                             3663 when "11010101010001",
                             3663 when "11010101010010",
                             3663 when "11010101010011",
                             3662 when "11010101010100",
                             3662 when "11010101010101",
                             3662 when "11010101010110",
                             3662 when "11010101010111",
                             3661 when "11010101011000",
                             3661 when "11010101011001",
                             3661 when "11010101011010",
                             3661 when "11010101011011",
                             3660 when "11010101011100",
                             3660 when "11010101011101",
                             3660 when "11010101011110",
                             3660 when "11010101011111",
                             3659 when "11010101100000",
                             3659 when "11010101100001",
                             3659 when "11010101100010",
                             3658 when "11010101100011",
                             3658 when "11010101100100",
                             3658 when "11010101100101",
                             3658 when "11010101100110",
                             3657 when "11010101100111",
                             3657 when "11010101101000",
                             3657 when "11010101101001",
                             3657 when "11010101101010",
                             3656 when "11010101101011",
                             3656 when "11010101101100",
                             3656 when "11010101101101",
                             3656 when "11010101101110",
                             3655 when "11010101101111",
                             3655 when "11010101110000",
                             3655 when "11010101110001",
                             3654 when "11010101110010",
                             3654 when "11010101110011",
                             3654 when "11010101110100",
                             3654 when "11010101110101",
                             3653 when "11010101110110",
                             3653 when "11010101110111",
                             3653 when "11010101111000",
                             3653 when "11010101111001",
                             3652 when "11010101111010",
                             3652 when "11010101111011",
                             3652 when "11010101111100",
                             3652 when "11010101111101",
                             3651 when "11010101111110",
                             3651 when "11010101111111",
                             3651 when "11010110000000",
                             3650 when "11010110000001",
                             3650 when "11010110000010",
                             3650 when "11010110000011",
                             3650 when "11010110000100",
                             3649 when "11010110000101",
                             3649 when "11010110000110",
                             3649 when "11010110000111",
                             3649 when "11010110001000",
                             3648 when "11010110001001",
                             3648 when "11010110001010",
                             3648 when "11010110001011",
                             3648 when "11010110001100",
                             3647 when "11010110001101",
                             3647 when "11010110001110",
                             3647 when "11010110001111",
                             3646 when "11010110010000",
                             3646 when "11010110010001",
                             3646 when "11010110010010",
                             3646 when "11010110010011",
                             3645 when "11010110010100",
                             3645 when "11010110010101",
                             3645 when "11010110010110",
                             3645 when "11010110010111",
                             3644 when "11010110011000",
                             3644 when "11010110011001",
                             3644 when "11010110011010",
                             3644 when "11010110011011",
                             3643 when "11010110011100",
                             3643 when "11010110011101",
                             3643 when "11010110011110",
                             3642 when "11010110011111",
                             3642 when "11010110100000",
                             3642 when "11010110100001",
                             3642 when "11010110100010",
                             3641 when "11010110100011",
                             3641 when "11010110100100",
                             3641 when "11010110100101",
                             3641 when "11010110100110",
                             3640 when "11010110100111",
                             3640 when "11010110101000",
                             3640 when "11010110101001",
                             3640 when "11010110101010",
                             3639 when "11010110101011",
                             3639 when "11010110101100",
                             3639 when "11010110101101",
                             3638 when "11010110101110",
                             3638 when "11010110101111",
                             3638 when "11010110110000",
                             3638 when "11010110110001",
                             3637 when "11010110110010",
                             3637 when "11010110110011",
                             3637 when "11010110110100",
                             3637 when "11010110110101",
                             3636 when "11010110110110",
                             3636 when "11010110110111",
                             3636 when "11010110111000",
                             3636 when "11010110111001",
                             3635 when "11010110111010",
                             3635 when "11010110111011",
                             3635 when "11010110111100",
                             3635 when "11010110111101",
                             3634 when "11010110111110",
                             3634 when "11010110111111",
                             3634 when "11010111000000",
                             3633 when "11010111000001",
                             3633 when "11010111000010",
                             3633 when "11010111000011",
                             3633 when "11010111000100",
                             3632 when "11010111000101",
                             3632 when "11010111000110",
                             3632 when "11010111000111",
                             3632 when "11010111001000",
                             3631 when "11010111001001",
                             3631 when "11010111001010",
                             3631 when "11010111001011",
                             3631 when "11010111001100",
                             3630 when "11010111001101",
                             3630 when "11010111001110",
                             3630 when "11010111001111",
                             3630 when "11010111010000",
                             3629 when "11010111010001",
                             3629 when "11010111010010",
                             3629 when "11010111010011",
                             3628 when "11010111010100",
                             3628 when "11010111010101",
                             3628 when "11010111010110",
                             3628 when "11010111010111",
                             3627 when "11010111011000",
                             3627 when "11010111011001",
                             3627 when "11010111011010",
                             3627 when "11010111011011",
                             3626 when "11010111011100",
                             3626 when "11010111011101",
                             3626 when "11010111011110",
                             3626 when "11010111011111",
                             3625 when "11010111100000",
                             3625 when "11010111100001",
                             3625 when "11010111100010",
                             3625 when "11010111100011",
                             3624 when "11010111100100",
                             3624 when "11010111100101",
                             3624 when "11010111100110",
                             3623 when "11010111100111",
                             3623 when "11010111101000",
                             3623 when "11010111101001",
                             3623 when "11010111101010",
                             3622 when "11010111101011",
                             3622 when "11010111101100",
                             3622 when "11010111101101",
                             3622 when "11010111101110",
                             3621 when "11010111101111",
                             3621 when "11010111110000",
                             3621 when "11010111110001",
                             3621 when "11010111110010",
                             3620 when "11010111110011",
                             3620 when "11010111110100",
                             3620 when "11010111110101",
                             3620 when "11010111110110",
                             3619 when "11010111110111",
                             3619 when "11010111111000",
                             3619 when "11010111111001",
                             3618 when "11010111111010",
                             3618 when "11010111111011",
                             3618 when "11010111111100",
                             3618 when "11010111111101",
                             3617 when "11010111111110",
                             3617 when "11010111111111",
                             3617 when "11011000000000",
                             3617 when "11011000000001",
                             3616 when "11011000000010",
                             3616 when "11011000000011",
                             3616 when "11011000000100",
                             3616 when "11011000000101",
                             3615 when "11011000000110",
                             3615 when "11011000000111",
                             3615 when "11011000001000",
                             3615 when "11011000001001",
                             3614 when "11011000001010",
                             3614 when "11011000001011",
                             3614 when "11011000001100",
                             3614 when "11011000001101",
                             3613 when "11011000001110",
                             3613 when "11011000001111",
                             3613 when "11011000010000",
                             3612 when "11011000010001",
                             3612 when "11011000010010",
                             3612 when "11011000010011",
                             3612 when "11011000010100",
                             3611 when "11011000010101",
                             3611 when "11011000010110",
                             3611 when "11011000010111",
                             3611 when "11011000011000",
                             3610 when "11011000011001",
                             3610 when "11011000011010",
                             3610 when "11011000011011",
                             3610 when "11011000011100",
                             3609 when "11011000011101",
                             3609 when "11011000011110",
                             3609 when "11011000011111",
                             3609 when "11011000100000",
                             3608 when "11011000100001",
                             3608 when "11011000100010",
                             3608 when "11011000100011",
                             3608 when "11011000100100",
                             3607 when "11011000100101",
                             3607 when "11011000100110",
                             3607 when "11011000100111",
                             3606 when "11011000101000",
                             3606 when "11011000101001",
                             3606 when "11011000101010",
                             3606 when "11011000101011",
                             3605 when "11011000101100",
                             3605 when "11011000101101",
                             3605 when "11011000101110",
                             3605 when "11011000101111",
                             3604 when "11011000110000",
                             3604 when "11011000110001",
                             3604 when "11011000110010",
                             3604 when "11011000110011",
                             3603 when "11011000110100",
                             3603 when "11011000110101",
                             3603 when "11011000110110",
                             3603 when "11011000110111",
                             3602 when "11011000111000",
                             3602 when "11011000111001",
                             3602 when "11011000111010",
                             3602 when "11011000111011",
                             3601 when "11011000111100",
                             3601 when "11011000111101",
                             3601 when "11011000111110",
                             3600 when "11011000111111",
                             3600 when "11011001000000",
                             3600 when "11011001000001",
                             3600 when "11011001000010",
                             3599 when "11011001000011",
                             3599 when "11011001000100",
                             3599 when "11011001000101",
                             3599 when "11011001000110",
                             3598 when "11011001000111",
                             3598 when "11011001001000",
                             3598 when "11011001001001",
                             3598 when "11011001001010",
                             3597 when "11011001001011",
                             3597 when "11011001001100",
                             3597 when "11011001001101",
                             3597 when "11011001001110",
                             3596 when "11011001001111",
                             3596 when "11011001010000",
                             3596 when "11011001010001",
                             3596 when "11011001010010",
                             3595 when "11011001010011",
                             3595 when "11011001010100",
                             3595 when "11011001010101",
                             3595 when "11011001010110",
                             3594 when "11011001010111",
                             3594 when "11011001011000",
                             3594 when "11011001011001",
                             3594 when "11011001011010",
                             3593 when "11011001011011",
                             3593 when "11011001011100",
                             3593 when "11011001011101",
                             3592 when "11011001011110",
                             3592 when "11011001011111",
                             3592 when "11011001100000",
                             3592 when "11011001100001",
                             3591 when "11011001100010",
                             3591 when "11011001100011",
                             3591 when "11011001100100",
                             3591 when "11011001100101",
                             3590 when "11011001100110",
                             3590 when "11011001100111",
                             3590 when "11011001101000",
                             3590 when "11011001101001",
                             3589 when "11011001101010",
                             3589 when "11011001101011",
                             3589 when "11011001101100",
                             3589 when "11011001101101",
                             3588 when "11011001101110",
                             3588 when "11011001101111",
                             3588 when "11011001110000",
                             3588 when "11011001110001",
                             3587 when "11011001110010",
                             3587 when "11011001110011",
                             3587 when "11011001110100",
                             3587 when "11011001110101",
                             3586 when "11011001110110",
                             3586 when "11011001110111",
                             3586 when "11011001111000",
                             3586 when "11011001111001",
                             3585 when "11011001111010",
                             3585 when "11011001111011",
                             3585 when "11011001111100",
                             3584 when "11011001111101",
                             3584 when "11011001111110",
                             3584 when "11011001111111",
                             3584 when "11011010000000",
                             3583 when "11011010000001",
                             3583 when "11011010000010",
                             3583 when "11011010000011",
                             3583 when "11011010000100",
                             3582 when "11011010000101",
                             3582 when "11011010000110",
                             3582 when "11011010000111",
                             3582 when "11011010001000",
                             3581 when "11011010001001",
                             3581 when "11011010001010",
                             3581 when "11011010001011",
                             3581 when "11011010001100",
                             3580 when "11011010001101",
                             3580 when "11011010001110",
                             3580 when "11011010001111",
                             3580 when "11011010010000",
                             3579 when "11011010010001",
                             3579 when "11011010010010",
                             3579 when "11011010010011",
                             3579 when "11011010010100",
                             3578 when "11011010010101",
                             3578 when "11011010010110",
                             3578 when "11011010010111",
                             3578 when "11011010011000",
                             3577 when "11011010011001",
                             3577 when "11011010011010",
                             3577 when "11011010011011",
                             3577 when "11011010011100",
                             3576 when "11011010011101",
                             3576 when "11011010011110",
                             3576 when "11011010011111",
                             3576 when "11011010100000",
                             3575 when "11011010100001",
                             3575 when "11011010100010",
                             3575 when "11011010100011",
                             3574 when "11011010100100",
                             3574 when "11011010100101",
                             3574 when "11011010100110",
                             3574 when "11011010100111",
                             3573 when "11011010101000",
                             3573 when "11011010101001",
                             3573 when "11011010101010",
                             3573 when "11011010101011",
                             3572 when "11011010101100",
                             3572 when "11011010101101",
                             3572 when "11011010101110",
                             3572 when "11011010101111",
                             3571 when "11011010110000",
                             3571 when "11011010110001",
                             3571 when "11011010110010",
                             3571 when "11011010110011",
                             3570 when "11011010110100",
                             3570 when "11011010110101",
                             3570 when "11011010110110",
                             3570 when "11011010110111",
                             3569 when "11011010111000",
                             3569 when "11011010111001",
                             3569 when "11011010111010",
                             3569 when "11011010111011",
                             3568 when "11011010111100",
                             3568 when "11011010111101",
                             3568 when "11011010111110",
                             3568 when "11011010111111",
                             3567 when "11011011000000",
                             3567 when "11011011000001",
                             3567 when "11011011000010",
                             3567 when "11011011000011",
                             3566 when "11011011000100",
                             3566 when "11011011000101",
                             3566 when "11011011000110",
                             3566 when "11011011000111",
                             3565 when "11011011001000",
                             3565 when "11011011001001",
                             3565 when "11011011001010",
                             3565 when "11011011001011",
                             3564 when "11011011001100",
                             3564 when "11011011001101",
                             3564 when "11011011001110",
                             3564 when "11011011001111",
                             3563 when "11011011010000",
                             3563 when "11011011010001",
                             3563 when "11011011010010",
                             3563 when "11011011010011",
                             3562 when "11011011010100",
                             3562 when "11011011010101",
                             3562 when "11011011010110",
                             3562 when "11011011010111",
                             3561 when "11011011011000",
                             3561 when "11011011011001",
                             3561 when "11011011011010",
                             3560 when "11011011011011",
                             3560 when "11011011011100",
                             3560 when "11011011011101",
                             3560 when "11011011011110",
                             3559 when "11011011011111",
                             3559 when "11011011100000",
                             3559 when "11011011100001",
                             3559 when "11011011100010",
                             3558 when "11011011100011",
                             3558 when "11011011100100",
                             3558 when "11011011100101",
                             3558 when "11011011100110",
                             3557 when "11011011100111",
                             3557 when "11011011101000",
                             3557 when "11011011101001",
                             3557 when "11011011101010",
                             3556 when "11011011101011",
                             3556 when "11011011101100",
                             3556 when "11011011101101",
                             3556 when "11011011101110",
                             3555 when "11011011101111",
                             3555 when "11011011110000",
                             3555 when "11011011110001",
                             3555 when "11011011110010",
                             3554 when "11011011110011",
                             3554 when "11011011110100",
                             3554 when "11011011110101",
                             3554 when "11011011110110",
                             3553 when "11011011110111",
                             3553 when "11011011111000",
                             3553 when "11011011111001",
                             3553 when "11011011111010",
                             3552 when "11011011111011",
                             3552 when "11011011111100",
                             3552 when "11011011111101",
                             3552 when "11011011111110",
                             3551 when "11011011111111",
                             3551 when "11011100000000",
                             3551 when "11011100000001",
                             3551 when "11011100000010",
                             3550 when "11011100000011",
                             3550 when "11011100000100",
                             3550 when "11011100000101",
                             3550 when "11011100000110",
                             3549 when "11011100000111",
                             3549 when "11011100001000",
                             3549 when "11011100001001",
                             3549 when "11011100001010",
                             3548 when "11011100001011",
                             3548 when "11011100001100",
                             3548 when "11011100001101",
                             3548 when "11011100001110",
                             3547 when "11011100001111",
                             3547 when "11011100010000",
                             3547 when "11011100010001",
                             3547 when "11011100010010",
                             3546 when "11011100010011",
                             3546 when "11011100010100",
                             3546 when "11011100010101",
                             3546 when "11011100010110",
                             3545 when "11011100010111",
                             3545 when "11011100011000",
                             3545 when "11011100011001",
                             3545 when "11011100011010",
                             3544 when "11011100011011",
                             3544 when "11011100011100",
                             3544 when "11011100011101",
                             3544 when "11011100011110",
                             3543 when "11011100011111",
                             3543 when "11011100100000",
                             3543 when "11011100100001",
                             3543 when "11011100100010",
                             3542 when "11011100100011",
                             3542 when "11011100100100",
                             3542 when "11011100100101",
                             3542 when "11011100100110",
                             3541 when "11011100100111",
                             3541 when "11011100101000",
                             3541 when "11011100101001",
                             3541 when "11011100101010",
                             3540 when "11011100101011",
                             3540 when "11011100101100",
                             3540 when "11011100101101",
                             3540 when "11011100101110",
                             3539 when "11011100101111",
                             3539 when "11011100110000",
                             3539 when "11011100110001",
                             3539 when "11011100110010",
                             3538 when "11011100110011",
                             3538 when "11011100110100",
                             3538 when "11011100110101",
                             3538 when "11011100110110",
                             3537 when "11011100110111",
                             3537 when "11011100111000",
                             3537 when "11011100111001",
                             3537 when "11011100111010",
                             3536 when "11011100111011",
                             3536 when "11011100111100",
                             3536 when "11011100111101",
                             3536 when "11011100111110",
                             3535 when "11011100111111",
                             3535 when "11011101000000",
                             3535 when "11011101000001",
                             3535 when "11011101000010",
                             3534 when "11011101000011",
                             3534 when "11011101000100",
                             3534 when "11011101000101",
                             3534 when "11011101000110",
                             3533 when "11011101000111",
                             3533 when "11011101001000",
                             3533 when "11011101001001",
                             3533 when "11011101001010",
                             3532 when "11011101001011",
                             3532 when "11011101001100",
                             3532 when "11011101001101",
                             3532 when "11011101001110",
                             3531 when "11011101001111",
                             3531 when "11011101010000",
                             3531 when "11011101010001",
                             3531 when "11011101010010",
                             3530 when "11011101010011",
                             3530 when "11011101010100",
                             3530 when "11011101010101",
                             3530 when "11011101010110",
                             3529 when "11011101010111",
                             3529 when "11011101011000",
                             3529 when "11011101011001",
                             3529 when "11011101011010",
                             3528 when "11011101011011",
                             3528 when "11011101011100",
                             3528 when "11011101011101",
                             3528 when "11011101011110",
                             3527 when "11011101011111",
                             3527 when "11011101100000",
                             3527 when "11011101100001",
                             3527 when "11011101100010",
                             3526 when "11011101100011",
                             3526 when "11011101100100",
                             3526 when "11011101100101",
                             3526 when "11011101100110",
                             3525 when "11011101100111",
                             3525 when "11011101101000",
                             3525 when "11011101101001",
                             3525 when "11011101101010",
                             3524 when "11011101101011",
                             3524 when "11011101101100",
                             3524 when "11011101101101",
                             3524 when "11011101101110",
                             3523 when "11011101101111",
                             3523 when "11011101110000",
                             3523 when "11011101110001",
                             3523 when "11011101110010",
                             3522 when "11011101110011",
                             3522 when "11011101110100",
                             3522 when "11011101110101",
                             3522 when "11011101110110",
                             3521 when "11011101110111",
                             3521 when "11011101111000",
                             3521 when "11011101111001",
                             3521 when "11011101111010",
                             3520 when "11011101111011",
                             3520 when "11011101111100",
                             3520 when "11011101111101",
                             3520 when "11011101111110",
                             3519 when "11011101111111",
                             3519 when "11011110000000",
                             3519 when "11011110000001",
                             3519 when "11011110000010",
                             3518 when "11011110000011",
                             3518 when "11011110000100",
                             3518 when "11011110000101",
                             3518 when "11011110000110",
                             3517 when "11011110000111",
                             3517 when "11011110001000",
                             3517 when "11011110001001",
                             3517 when "11011110001010",
                             3516 when "11011110001011",
                             3516 when "11011110001100",
                             3516 when "11011110001101",
                             3516 when "11011110001110",
                             3515 when "11011110001111",
                             3515 when "11011110010000",
                             3515 when "11011110010001",
                             3515 when "11011110010010",
                             3514 when "11011110010011",
                             3514 when "11011110010100",
                             3514 when "11011110010101",
                             3514 when "11011110010110",
                             3513 when "11011110010111",
                             3513 when "11011110011000",
                             3513 when "11011110011001",
                             3513 when "11011110011010",
                             3512 when "11011110011011",
                             3512 when "11011110011100",
                             3512 when "11011110011101",
                             3512 when "11011110011110",
                             3511 when "11011110011111",
                             3511 when "11011110100000",
                             3511 when "11011110100001",
                             3511 when "11011110100010",
                             3510 when "11011110100011",
                             3510 when "11011110100100",
                             3510 when "11011110100101",
                             3510 when "11011110100110",
                             3510 when "11011110100111",
                             3509 when "11011110101000",
                             3509 when "11011110101001",
                             3509 when "11011110101010",
                             3509 when "11011110101011",
                             3508 when "11011110101100",
                             3508 when "11011110101101",
                             3508 when "11011110101110",
                             3508 when "11011110101111",
                             3507 when "11011110110000",
                             3507 when "11011110110001",
                             3507 when "11011110110010",
                             3507 when "11011110110011",
                             3506 when "11011110110100",
                             3506 when "11011110110101",
                             3506 when "11011110110110",
                             3506 when "11011110110111",
                             3505 when "11011110111000",
                             3505 when "11011110111001",
                             3505 when "11011110111010",
                             3505 when "11011110111011",
                             3504 when "11011110111100",
                             3504 when "11011110111101",
                             3504 when "11011110111110",
                             3504 when "11011110111111",
                             3503 when "11011111000000",
                             3503 when "11011111000001",
                             3503 when "11011111000010",
                             3503 when "11011111000011",
                             3502 when "11011111000100",
                             3502 when "11011111000101",
                             3502 when "11011111000110",
                             3502 when "11011111000111",
                             3501 when "11011111001000",
                             3501 when "11011111001001",
                             3501 when "11011111001010",
                             3501 when "11011111001011",
                             3500 when "11011111001100",
                             3500 when "11011111001101",
                             3500 when "11011111001110",
                             3500 when "11011111001111",
                             3499 when "11011111010000",
                             3499 when "11011111010001",
                             3499 when "11011111010010",
                             3499 when "11011111010011",
                             3498 when "11011111010100",
                             3498 when "11011111010101",
                             3498 when "11011111010110",
                             3498 when "11011111010111",
                             3497 when "11011111011000",
                             3497 when "11011111011001",
                             3497 when "11011111011010",
                             3497 when "11011111011011",
                             3497 when "11011111011100",
                             3496 when "11011111011101",
                             3496 when "11011111011110",
                             3496 when "11011111011111",
                             3496 when "11011111100000",
                             3495 when "11011111100001",
                             3495 when "11011111100010",
                             3495 when "11011111100011",
                             3495 when "11011111100100",
                             3494 when "11011111100101",
                             3494 when "11011111100110",
                             3494 when "11011111100111",
                             3494 when "11011111101000",
                             3493 when "11011111101001",
                             3493 when "11011111101010",
                             3493 when "11011111101011",
                             3493 when "11011111101100",
                             3492 when "11011111101101",
                             3492 when "11011111101110",
                             3492 when "11011111101111",
                             3492 when "11011111110000",
                             3491 when "11011111110001",
                             3491 when "11011111110010",
                             3491 when "11011111110011",
                             3491 when "11011111110100",
                             3490 when "11011111110101",
                             3490 when "11011111110110",
                             3490 when "11011111110111",
                             3490 when "11011111111000",
                             3489 when "11011111111001",
                             3489 when "11011111111010",
                             3489 when "11011111111011",
                             3489 when "11011111111100",
                             3488 when "11011111111101",
                             3488 when "11011111111110",
                             3488 when "11011111111111",
                             3488 when "11100000000000",
                             3487 when "11100000000001",
                             3487 when "11100000000010",
                             3487 when "11100000000011",
                             3487 when "11100000000100",
                             3487 when "11100000000101",
                             3486 when "11100000000110",
                             3486 when "11100000000111",
                             3486 when "11100000001000",
                             3486 when "11100000001001",
                             3485 when "11100000001010",
                             3485 when "11100000001011",
                             3485 when "11100000001100",
                             3485 when "11100000001101",
                             3484 when "11100000001110",
                             3484 when "11100000001111",
                             3484 when "11100000010000",
                             3484 when "11100000010001",
                             3483 when "11100000010010",
                             3483 when "11100000010011",
                             3483 when "11100000010100",
                             3483 when "11100000010101",
                             3482 when "11100000010110",
                             3482 when "11100000010111",
                             3482 when "11100000011000",
                             3482 when "11100000011001",
                             3481 when "11100000011010",
                             3481 when "11100000011011",
                             3481 when "11100000011100",
                             3481 when "11100000011101",
                             3480 when "11100000011110",
                             3480 when "11100000011111",
                             3480 when "11100000100000",
                             3480 when "11100000100001",
                             3479 when "11100000100010",
                             3479 when "11100000100011",
                             3479 when "11100000100100",
                             3479 when "11100000100101",
                             3479 when "11100000100110",
                             3478 when "11100000100111",
                             3478 when "11100000101000",
                             3478 when "11100000101001",
                             3478 when "11100000101010",
                             3477 when "11100000101011",
                             3477 when "11100000101100",
                             3477 when "11100000101101",
                             3477 when "11100000101110",
                             3476 when "11100000101111",
                             3476 when "11100000110000",
                             3476 when "11100000110001",
                             3476 when "11100000110010",
                             3475 when "11100000110011",
                             3475 when "11100000110100",
                             3475 when "11100000110101",
                             3475 when "11100000110110",
                             3474 when "11100000110111",
                             3474 when "11100000111000",
                             3474 when "11100000111001",
                             3474 when "11100000111010",
                             3473 when "11100000111011",
                             3473 when "11100000111100",
                             3473 when "11100000111101",
                             3473 when "11100000111110",
                             3472 when "11100000111111",
                             3472 when "11100001000000",
                             3472 when "11100001000001",
                             3472 when "11100001000010",
                             3471 when "11100001000011",
                             3471 when "11100001000100",
                             3471 when "11100001000101",
                             3471 when "11100001000110",
                             3471 when "11100001000111",
                             3470 when "11100001001000",
                             3470 when "11100001001001",
                             3470 when "11100001001010",
                             3470 when "11100001001011",
                             3469 when "11100001001100",
                             3469 when "11100001001101",
                             3469 when "11100001001110",
                             3469 when "11100001001111",
                             3468 when "11100001010000",
                             3468 when "11100001010001",
                             3468 when "11100001010010",
                             3468 when "11100001010011",
                             3467 when "11100001010100",
                             3467 when "11100001010101",
                             3467 when "11100001010110",
                             3467 when "11100001010111",
                             3466 when "11100001011000",
                             3466 when "11100001011001",
                             3466 when "11100001011010",
                             3466 when "11100001011011",
                             3465 when "11100001011100",
                             3465 when "11100001011101",
                             3465 when "11100001011110",
                             3465 when "11100001011111",
                             3465 when "11100001100000",
                             3464 when "11100001100001",
                             3464 when "11100001100010",
                             3464 when "11100001100011",
                             3464 when "11100001100100",
                             3463 when "11100001100101",
                             3463 when "11100001100110",
                             3463 when "11100001100111",
                             3463 when "11100001101000",
                             3462 when "11100001101001",
                             3462 when "11100001101010",
                             3462 when "11100001101011",
                             3462 when "11100001101100",
                             3461 when "11100001101101",
                             3461 when "11100001101110",
                             3461 when "11100001101111",
                             3461 when "11100001110000",
                             3460 when "11100001110001",
                             3460 when "11100001110010",
                             3460 when "11100001110011",
                             3460 when "11100001110100",
                             3459 when "11100001110101",
                             3459 when "11100001110110",
                             3459 when "11100001110111",
                             3459 when "11100001111000",
                             3459 when "11100001111001",
                             3458 when "11100001111010",
                             3458 when "11100001111011",
                             3458 when "11100001111100",
                             3458 when "11100001111101",
                             3457 when "11100001111110",
                             3457 when "11100001111111",
                             3457 when "11100010000000",
                             3457 when "11100010000001",
                             3456 when "11100010000010",
                             3456 when "11100010000011",
                             3456 when "11100010000100",
                             3456 when "11100010000101",
                             3455 when "11100010000110",
                             3455 when "11100010000111",
                             3455 when "11100010001000",
                             3455 when "11100010001001",
                             3454 when "11100010001010",
                             3454 when "11100010001011",
                             3454 when "11100010001100",
                             3454 when "11100010001101",
                             3454 when "11100010001110",
                             3453 when "11100010001111",
                             3453 when "11100010010000",
                             3453 when "11100010010001",
                             3453 when "11100010010010",
                             3452 when "11100010010011",
                             3452 when "11100010010100",
                             3452 when "11100010010101",
                             3452 when "11100010010110",
                             3451 when "11100010010111",
                             3451 when "11100010011000",
                             3451 when "11100010011001",
                             3451 when "11100010011010",
                             3450 when "11100010011011",
                             3450 when "11100010011100",
                             3450 when "11100010011101",
                             3450 when "11100010011110",
                             3449 when "11100010011111",
                             3449 when "11100010100000",
                             3449 when "11100010100001",
                             3449 when "11100010100010",
                             3449 when "11100010100011",
                             3448 when "11100010100100",
                             3448 when "11100010100101",
                             3448 when "11100010100110",
                             3448 when "11100010100111",
                             3447 when "11100010101000",
                             3447 when "11100010101001",
                             3447 when "11100010101010",
                             3447 when "11100010101011",
                             3446 when "11100010101100",
                             3446 when "11100010101101",
                             3446 when "11100010101110",
                             3446 when "11100010101111",
                             3445 when "11100010110000",
                             3445 when "11100010110001",
                             3445 when "11100010110010",
                             3445 when "11100010110011",
                             3444 when "11100010110100",
                             3444 when "11100010110101",
                             3444 when "11100010110110",
                             3444 when "11100010110111",
                             3444 when "11100010111000",
                             3443 when "11100010111001",
                             3443 when "11100010111010",
                             3443 when "11100010111011",
                             3443 when "11100010111100",
                             3442 when "11100010111101",
                             3442 when "11100010111110",
                             3442 when "11100010111111",
                             3442 when "11100011000000",
                             3441 when "11100011000001",
                             3441 when "11100011000010",
                             3441 when "11100011000011",
                             3441 when "11100011000100",
                             3440 when "11100011000101",
                             3440 when "11100011000110",
                             3440 when "11100011000111",
                             3440 when "11100011001000",
                             3439 when "11100011001001",
                             3439 when "11100011001010",
                             3439 when "11100011001011",
                             3439 when "11100011001100",
                             3439 when "11100011001101",
                             3438 when "11100011001110",
                             3438 when "11100011001111",
                             3438 when "11100011010000",
                             3438 when "11100011010001",
                             3437 when "11100011010010",
                             3437 when "11100011010011",
                             3437 when "11100011010100",
                             3437 when "11100011010101",
                             3436 when "11100011010110",
                             3436 when "11100011010111",
                             3436 when "11100011011000",
                             3436 when "11100011011001",
                             3435 when "11100011011010",
                             3435 when "11100011011011",
                             3435 when "11100011011100",
                             3435 when "11100011011101",
                             3435 when "11100011011110",
                             3434 when "11100011011111",
                             3434 when "11100011100000",
                             3434 when "11100011100001",
                             3434 when "11100011100010",
                             3433 when "11100011100011",
                             3433 when "11100011100100",
                             3433 when "11100011100101",
                             3433 when "11100011100110",
                             3432 when "11100011100111",
                             3432 when "11100011101000",
                             3432 when "11100011101001",
                             3432 when "11100011101010",
                             3431 when "11100011101011",
                             3431 when "11100011101100",
                             3431 when "11100011101101",
                             3431 when "11100011101110",
                             3431 when "11100011101111",
                             3430 when "11100011110000",
                             3430 when "11100011110001",
                             3430 when "11100011110010",
                             3430 when "11100011110011",
                             3429 when "11100011110100",
                             3429 when "11100011110101",
                             3429 when "11100011110110",
                             3429 when "11100011110111",
                             3428 when "11100011111000",
                             3428 when "11100011111001",
                             3428 when "11100011111010",
                             3428 when "11100011111011",
                             3427 when "11100011111100",
                             3427 when "11100011111101",
                             3427 when "11100011111110",
                             3427 when "11100011111111",
                             3427 when "11100100000000",
                             3426 when "11100100000001",
                             3426 when "11100100000010",
                             3426 when "11100100000011",
                             3426 when "11100100000100",
                             3425 when "11100100000101",
                             3425 when "11100100000110",
                             3425 when "11100100000111",
                             3425 when "11100100001000",
                             3424 when "11100100001001",
                             3424 when "11100100001010",
                             3424 when "11100100001011",
                             3424 when "11100100001100",
                             3423 when "11100100001101",
                             3423 when "11100100001110",
                             3423 when "11100100001111",
                             3423 when "11100100010000",
                             3423 when "11100100010001",
                             3422 when "11100100010010",
                             3422 when "11100100010011",
                             3422 when "11100100010100",
                             3422 when "11100100010101",
                             3421 when "11100100010110",
                             3421 when "11100100010111",
                             3421 when "11100100011000",
                             3421 when "11100100011001",
                             3420 when "11100100011010",
                             3420 when "11100100011011",
                             3420 when "11100100011100",
                             3420 when "11100100011101",
                             3420 when "11100100011110",
                             3419 when "11100100011111",
                             3419 when "11100100100000",
                             3419 when "11100100100001",
                             3419 when "11100100100010",
                             3418 when "11100100100011",
                             3418 when "11100100100100",
                             3418 when "11100100100101",
                             3418 when "11100100100110",
                             3417 when "11100100100111",
                             3417 when "11100100101000",
                             3417 when "11100100101001",
                             3417 when "11100100101010",
                             3416 when "11100100101011",
                             3416 when "11100100101100",
                             3416 when "11100100101101",
                             3416 when "11100100101110",
                             3416 when "11100100101111",
                             3415 when "11100100110000",
                             3415 when "11100100110001",
                             3415 when "11100100110010",
                             3415 when "11100100110011",
                             3414 when "11100100110100",
                             3414 when "11100100110101",
                             3414 when "11100100110110",
                             3414 when "11100100110111",
                             3413 when "11100100111000",
                             3413 when "11100100111001",
                             3413 when "11100100111010",
                             3413 when "11100100111011",
                             3413 when "11100100111100",
                             3412 when "11100100111101",
                             3412 when "11100100111110",
                             3412 when "11100100111111",
                             3412 when "11100101000000",
                             3411 when "11100101000001",
                             3411 when "11100101000010",
                             3411 when "11100101000011",
                             3411 when "11100101000100",
                             3410 when "11100101000101",
                             3410 when "11100101000110",
                             3410 when "11100101000111",
                             3410 when "11100101001000",
                             3409 when "11100101001001",
                             3409 when "11100101001010",
                             3409 when "11100101001011",
                             3409 when "11100101001100",
                             3409 when "11100101001101",
                             3408 when "11100101001110",
                             3408 when "11100101001111",
                             3408 when "11100101010000",
                             3408 when "11100101010001",
                             3407 when "11100101010010",
                             3407 when "11100101010011",
                             3407 when "11100101010100",
                             3407 when "11100101010101",
                             3406 when "11100101010110",
                             3406 when "11100101010111",
                             3406 when "11100101011000",
                             3406 when "11100101011001",
                             3406 when "11100101011010",
                             3405 when "11100101011011",
                             3405 when "11100101011100",
                             3405 when "11100101011101",
                             3405 when "11100101011110",
                             3404 when "11100101011111",
                             3404 when "11100101100000",
                             3404 when "11100101100001",
                             3404 when "11100101100010",
                             3403 when "11100101100011",
                             3403 when "11100101100100",
                             3403 when "11100101100101",
                             3403 when "11100101100110",
                             3403 when "11100101100111",
                             3402 when "11100101101000",
                             3402 when "11100101101001",
                             3402 when "11100101101010",
                             3402 when "11100101101011",
                             3401 when "11100101101100",
                             3401 when "11100101101101",
                             3401 when "11100101101110",
                             3401 when "11100101101111",
                             3400 when "11100101110000",
                             3400 when "11100101110001",
                             3400 when "11100101110010",
                             3400 when "11100101110011",
                             3400 when "11100101110100",
                             3399 when "11100101110101",
                             3399 when "11100101110110",
                             3399 when "11100101110111",
                             3399 when "11100101111000",
                             3398 when "11100101111001",
                             3398 when "11100101111010",
                             3398 when "11100101111011",
                             3398 when "11100101111100",
                             3397 when "11100101111101",
                             3397 when "11100101111110",
                             3397 when "11100101111111",
                             3397 when "11100110000000",
                             3397 when "11100110000001",
                             3396 when "11100110000010",
                             3396 when "11100110000011",
                             3396 when "11100110000100",
                             3396 when "11100110000101",
                             3395 when "11100110000110",
                             3395 when "11100110000111",
                             3395 when "11100110001000",
                             3395 when "11100110001001",
                             3394 when "11100110001010",
                             3394 when "11100110001011",
                             3394 when "11100110001100",
                             3394 when "11100110001101",
                             3394 when "11100110001110",
                             3393 when "11100110001111",
                             3393 when "11100110010000",
                             3393 when "11100110010001",
                             3393 when "11100110010010",
                             3392 when "11100110010011",
                             3392 when "11100110010100",
                             3392 when "11100110010101",
                             3392 when "11100110010110",
                             3391 when "11100110010111",
                             3391 when "11100110011000",
                             3391 when "11100110011001",
                             3391 when "11100110011010",
                             3391 when "11100110011011",
                             3390 when "11100110011100",
                             3390 when "11100110011101",
                             3390 when "11100110011110",
                             3390 when "11100110011111",
                             3389 when "11100110100000",
                             3389 when "11100110100001",
                             3389 when "11100110100010",
                             3389 when "11100110100011",
                             3388 when "11100110100100",
                             3388 when "11100110100101",
                             3388 when "11100110100110",
                             3388 when "11100110100111",
                             3388 when "11100110101000",
                             3387 when "11100110101001",
                             3387 when "11100110101010",
                             3387 when "11100110101011",
                             3387 when "11100110101100",
                             3386 when "11100110101101",
                             3386 when "11100110101110",
                             3386 when "11100110101111",
                             3386 when "11100110110000",
                             3385 when "11100110110001",
                             3385 when "11100110110010",
                             3385 when "11100110110011",
                             3385 when "11100110110100",
                             3385 when "11100110110101",
                             3384 when "11100110110110",
                             3384 when "11100110110111",
                             3384 when "11100110111000",
                             3384 when "11100110111001",
                             3383 when "11100110111010",
                             3383 when "11100110111011",
                             3383 when "11100110111100",
                             3383 when "11100110111101",
                             3382 when "11100110111110",
                             3382 when "11100110111111",
                             3382 when "11100111000000",
                             3382 when "11100111000001",
                             3382 when "11100111000010",
                             3381 when "11100111000011",
                             3381 when "11100111000100",
                             3381 when "11100111000101",
                             3381 when "11100111000110",
                             3380 when "11100111000111",
                             3380 when "11100111001000",
                             3380 when "11100111001001",
                             3380 when "11100111001010",
                             3380 when "11100111001011",
                             3379 when "11100111001100",
                             3379 when "11100111001101",
                             3379 when "11100111001110",
                             3379 when "11100111001111",
                             3378 when "11100111010000",
                             3378 when "11100111010001",
                             3378 when "11100111010010",
                             3378 when "11100111010011",
                             3377 when "11100111010100",
                             3377 when "11100111010101",
                             3377 when "11100111010110",
                             3377 when "11100111010111",
                             3377 when "11100111011000",
                             3376 when "11100111011001",
                             3376 when "11100111011010",
                             3376 when "11100111011011",
                             3376 when "11100111011100",
                             3375 when "11100111011101",
                             3375 when "11100111011110",
                             3375 when "11100111011111",
                             3375 when "11100111100000",
                             3375 when "11100111100001",
                             3374 when "11100111100010",
                             3374 when "11100111100011",
                             3374 when "11100111100100",
                             3374 when "11100111100101",
                             3373 when "11100111100110",
                             3373 when "11100111100111",
                             3373 when "11100111101000",
                             3373 when "11100111101001",
                             3372 when "11100111101010",
                             3372 when "11100111101011",
                             3372 when "11100111101100",
                             3372 when "11100111101101",
                             3372 when "11100111101110",
                             3371 when "11100111101111",
                             3371 when "11100111110000",
                             3371 when "11100111110001",
                             3371 when "11100111110010",
                             3370 when "11100111110011",
                             3370 when "11100111110100",
                             3370 when "11100111110101",
                             3370 when "11100111110110",
                             3369 when "11100111110111",
                             3369 when "11100111111000",
                             3369 when "11100111111001",
                             3369 when "11100111111010",
                             3369 when "11100111111011",
                             3368 when "11100111111100",
                             3368 when "11100111111101",
                             3368 when "11100111111110",
                             3368 when "11100111111111",
                             3367 when "11101000000000",
                             3367 when "11101000000001",
                             3367 when "11101000000010",
                             3367 when "11101000000011",
                             3367 when "11101000000100",
                             3366 when "11101000000101",
                             3366 when "11101000000110",
                             3366 when "11101000000111",
                             3366 when "11101000001000",
                             3365 when "11101000001001",
                             3365 when "11101000001010",
                             3365 when "11101000001011",
                             3365 when "11101000001100",
                             3365 when "11101000001101",
                             3364 when "11101000001110",
                             3364 when "11101000001111",
                             3364 when "11101000010000",
                             3364 when "11101000010001",
                             3363 when "11101000010010",
                             3363 when "11101000010011",
                             3363 when "11101000010100",
                             3363 when "11101000010101",
                             3362 when "11101000010110",
                             3362 when "11101000010111",
                             3362 when "11101000011000",
                             3362 when "11101000011001",
                             3362 when "11101000011010",
                             3361 when "11101000011011",
                             3361 when "11101000011100",
                             3361 when "11101000011101",
                             3361 when "11101000011110",
                             3360 when "11101000011111",
                             3360 when "11101000100000",
                             3360 when "11101000100001",
                             3360 when "11101000100010",
                             3360 when "11101000100011",
                             3359 when "11101000100100",
                             3359 when "11101000100101",
                             3359 when "11101000100110",
                             3359 when "11101000100111",
                             3358 when "11101000101000",
                             3358 when "11101000101001",
                             3358 when "11101000101010",
                             3358 when "11101000101011",
                             3358 when "11101000101100",
                             3357 when "11101000101101",
                             3357 when "11101000101110",
                             3357 when "11101000101111",
                             3357 when "11101000110000",
                             3356 when "11101000110001",
                             3356 when "11101000110010",
                             3356 when "11101000110011",
                             3356 when "11101000110100",
                             3355 when "11101000110101",
                             3355 when "11101000110110",
                             3355 when "11101000110111",
                             3355 when "11101000111000",
                             3355 when "11101000111001",
                             3354 when "11101000111010",
                             3354 when "11101000111011",
                             3354 when "11101000111100",
                             3354 when "11101000111101",
                             3353 when "11101000111110",
                             3353 when "11101000111111",
                             3353 when "11101001000000",
                             3353 when "11101001000001",
                             3353 when "11101001000010",
                             3352 when "11101001000011",
                             3352 when "11101001000100",
                             3352 when "11101001000101",
                             3352 when "11101001000110",
                             3351 when "11101001000111",
                             3351 when "11101001001000",
                             3351 when "11101001001001",
                             3351 when "11101001001010",
                             3351 when "11101001001011",
                             3350 when "11101001001100",
                             3350 when "11101001001101",
                             3350 when "11101001001110",
                             3350 when "11101001001111",
                             3349 when "11101001010000",
                             3349 when "11101001010001",
                             3349 when "11101001010010",
                             3349 when "11101001010011",
                             3349 when "11101001010100",
                             3348 when "11101001010101",
                             3348 when "11101001010110",
                             3348 when "11101001010111",
                             3348 when "11101001011000",
                             3347 when "11101001011001",
                             3347 when "11101001011010",
                             3347 when "11101001011011",
                             3347 when "11101001011100",
                             3346 when "11101001011101",
                             3346 when "11101001011110",
                             3346 when "11101001011111",
                             3346 when "11101001100000",
                             3346 when "11101001100001",
                             3345 when "11101001100010",
                             3345 when "11101001100011",
                             3345 when "11101001100100",
                             3345 when "11101001100101",
                             3344 when "11101001100110",
                             3344 when "11101001100111",
                             3344 when "11101001101000",
                             3344 when "11101001101001",
                             3344 when "11101001101010",
                             3343 when "11101001101011",
                             3343 when "11101001101100",
                             3343 when "11101001101101",
                             3343 when "11101001101110",
                             3342 when "11101001101111",
                             3342 when "11101001110000",
                             3342 when "11101001110001",
                             3342 when "11101001110010",
                             3342 when "11101001110011",
                             3341 when "11101001110100",
                             3341 when "11101001110101",
                             3341 when "11101001110110",
                             3341 when "11101001110111",
                             3340 when "11101001111000",
                             3340 when "11101001111001",
                             3340 when "11101001111010",
                             3340 when "11101001111011",
                             3340 when "11101001111100",
                             3339 when "11101001111101",
                             3339 when "11101001111110",
                             3339 when "11101001111111",
                             3339 when "11101010000000",
                             3338 when "11101010000001",
                             3338 when "11101010000010",
                             3338 when "11101010000011",
                             3338 when "11101010000100",
                             3338 when "11101010000101",
                             3337 when "11101010000110",
                             3337 when "11101010000111",
                             3337 when "11101010001000",
                             3337 when "11101010001001",
                             3336 when "11101010001010",
                             3336 when "11101010001011",
                             3336 when "11101010001100",
                             3336 when "11101010001101",
                             3336 when "11101010001110",
                             3335 when "11101010001111",
                             3335 when "11101010010000",
                             3335 when "11101010010001",
                             3335 when "11101010010010",
                             3334 when "11101010010011",
                             3334 when "11101010010100",
                             3334 when "11101010010101",
                             3334 when "11101010010110",
                             3334 when "11101010010111",
                             3333 when "11101010011000",
                             3333 when "11101010011001",
                             3333 when "11101010011010",
                             3333 when "11101010011011",
                             3332 when "11101010011100",
                             3332 when "11101010011101",
                             3332 when "11101010011110",
                             3332 when "11101010011111",
                             3332 when "11101010100000",
                             3331 when "11101010100001",
                             3331 when "11101010100010",
                             3331 when "11101010100011",
                             3331 when "11101010100100",
                             3330 when "11101010100101",
                             3330 when "11101010100110",
                             3330 when "11101010100111",
                             3330 when "11101010101000",
                             3330 when "11101010101001",
                             3329 when "11101010101010",
                             3329 when "11101010101011",
                             3329 when "11101010101100",
                             3329 when "11101010101101",
                             3328 when "11101010101110",
                             3328 when "11101010101111",
                             3328 when "11101010110000",
                             3328 when "11101010110001",
                             3328 when "11101010110010",
                             3327 when "11101010110011",
                             3327 when "11101010110100",
                             3327 when "11101010110101",
                             3327 when "11101010110110",
                             3326 when "11101010110111",
                             3326 when "11101010111000",
                             3326 when "11101010111001",
                             3326 when "11101010111010",
                             3326 when "11101010111011",
                             3325 when "11101010111100",
                             3325 when "11101010111101",
                             3325 when "11101010111110",
                             3325 when "11101010111111",
                             3324 when "11101011000000",
                             3324 when "11101011000001",
                             3324 when "11101011000010",
                             3324 when "11101011000011",
                             3324 when "11101011000100",
                             3323 when "11101011000101",
                             3323 when "11101011000110",
                             3323 when "11101011000111",
                             3323 when "11101011001000",
                             3322 when "11101011001001",
                             3322 when "11101011001010",
                             3322 when "11101011001011",
                             3322 when "11101011001100",
                             3322 when "11101011001101",
                             3321 when "11101011001110",
                             3321 when "11101011001111",
                             3321 when "11101011010000",
                             3321 when "11101011010001",
                             3320 when "11101011010010",
                             3320 when "11101011010011",
                             3320 when "11101011010100",
                             3320 when "11101011010101",
                             3320 when "11101011010110",
                             3319 when "11101011010111",
                             3319 when "11101011011000",
                             3319 when "11101011011001",
                             3319 when "11101011011010",
                             3319 when "11101011011011",
                             3318 when "11101011011100",
                             3318 when "11101011011101",
                             3318 when "11101011011110",
                             3318 when "11101011011111",
                             3317 when "11101011100000",
                             3317 when "11101011100001",
                             3317 when "11101011100010",
                             3317 when "11101011100011",
                             3317 when "11101011100100",
                             3316 when "11101011100101",
                             3316 when "11101011100110",
                             3316 when "11101011100111",
                             3316 when "11101011101000",
                             3315 when "11101011101001",
                             3315 when "11101011101010",
                             3315 when "11101011101011",
                             3315 when "11101011101100",
                             3315 when "11101011101101",
                             3314 when "11101011101110",
                             3314 when "11101011101111",
                             3314 when "11101011110000",
                             3314 when "11101011110001",
                             3313 when "11101011110010",
                             3313 when "11101011110011",
                             3313 when "11101011110100",
                             3313 when "11101011110101",
                             3313 when "11101011110110",
                             3312 when "11101011110111",
                             3312 when "11101011111000",
                             3312 when "11101011111001",
                             3312 when "11101011111010",
                             3311 when "11101011111011",
                             3311 when "11101011111100",
                             3311 when "11101011111101",
                             3311 when "11101011111110",
                             3311 when "11101011111111",
                             3310 when "11101100000000",
                             3310 when "11101100000001",
                             3310 when "11101100000010",
                             3310 when "11101100000011",
                             3310 when "11101100000100",
                             3309 when "11101100000101",
                             3309 when "11101100000110",
                             3309 when "11101100000111",
                             3309 when "11101100001000",
                             3308 when "11101100001001",
                             3308 when "11101100001010",
                             3308 when "11101100001011",
                             3308 when "11101100001100",
                             3308 when "11101100001101",
                             3307 when "11101100001110",
                             3307 when "11101100001111",
                             3307 when "11101100010000",
                             3307 when "11101100010001",
                             3306 when "11101100010010",
                             3306 when "11101100010011",
                             3306 when "11101100010100",
                             3306 when "11101100010101",
                             3306 when "11101100010110",
                             3305 when "11101100010111",
                             3305 when "11101100011000",
                             3305 when "11101100011001",
                             3305 when "11101100011010",
                             3304 when "11101100011011",
                             3304 when "11101100011100",
                             3304 when "11101100011101",
                             3304 when "11101100011110",
                             3304 when "11101100011111",
                             3303 when "11101100100000",
                             3303 when "11101100100001",
                             3303 when "11101100100010",
                             3303 when "11101100100011",
                             3303 when "11101100100100",
                             3302 when "11101100100101",
                             3302 when "11101100100110",
                             3302 when "11101100100111",
                             3302 when "11101100101000",
                             3301 when "11101100101001",
                             3301 when "11101100101010",
                             3301 when "11101100101011",
                             3301 when "11101100101100",
                             3301 when "11101100101101",
                             3300 when "11101100101110",
                             3300 when "11101100101111",
                             3300 when "11101100110000",
                             3300 when "11101100110001",
                             3299 when "11101100110010",
                             3299 when "11101100110011",
                             3299 when "11101100110100",
                             3299 when "11101100110101",
                             3299 when "11101100110110",
                             3298 when "11101100110111",
                             3298 when "11101100111000",
                             3298 when "11101100111001",
                             3298 when "11101100111010",
                             3298 when "11101100111011",
                             3297 when "11101100111100",
                             3297 when "11101100111101",
                             3297 when "11101100111110",
                             3297 when "11101100111111",
                             3296 when "11101101000000",
                             3296 when "11101101000001",
                             3296 when "11101101000010",
                             3296 when "11101101000011",
                             3296 when "11101101000100",
                             3295 when "11101101000101",
                             3295 when "11101101000110",
                             3295 when "11101101000111",
                             3295 when "11101101001000",
                             3294 when "11101101001001",
                             3294 when "11101101001010",
                             3294 when "11101101001011",
                             3294 when "11101101001100",
                             3294 when "11101101001101",
                             3293 when "11101101001110",
                             3293 when "11101101001111",
                             3293 when "11101101010000",
                             3293 when "11101101010001",
                             3293 when "11101101010010",
                             3292 when "11101101010011",
                             3292 when "11101101010100",
                             3292 when "11101101010101",
                             3292 when "11101101010110",
                             3291 when "11101101010111",
                             3291 when "11101101011000",
                             3291 when "11101101011001",
                             3291 when "11101101011010",
                             3291 when "11101101011011",
                             3290 when "11101101011100",
                             3290 when "11101101011101",
                             3290 when "11101101011110",
                             3290 when "11101101011111",
                             3289 when "11101101100000",
                             3289 when "11101101100001",
                             3289 when "11101101100010",
                             3289 when "11101101100011",
                             3289 when "11101101100100",
                             3288 when "11101101100101",
                             3288 when "11101101100110",
                             3288 when "11101101100111",
                             3288 when "11101101101000",
                             3288 when "11101101101001",
                             3287 when "11101101101010",
                             3287 when "11101101101011",
                             3287 when "11101101101100",
                             3287 when "11101101101101",
                             3286 when "11101101101110",
                             3286 when "11101101101111",
                             3286 when "11101101110000",
                             3286 when "11101101110001",
                             3286 when "11101101110010",
                             3285 when "11101101110011",
                             3285 when "11101101110100",
                             3285 when "11101101110101",
                             3285 when "11101101110110",
                             3285 when "11101101110111",
                             3284 when "11101101111000",
                             3284 when "11101101111001",
                             3284 when "11101101111010",
                             3284 when "11101101111011",
                             3283 when "11101101111100",
                             3283 when "11101101111101",
                             3283 when "11101101111110",
                             3283 when "11101101111111",
                             3283 when "11101110000000",
                             3282 when "11101110000001",
                             3282 when "11101110000010",
                             3282 when "11101110000011",
                             3282 when "11101110000100",
                             3281 when "11101110000101",
                             3281 when "11101110000110",
                             3281 when "11101110000111",
                             3281 when "11101110001000",
                             3281 when "11101110001001",
                             3280 when "11101110001010",
                             3280 when "11101110001011",
                             3280 when "11101110001100",
                             3280 when "11101110001101",
                             3280 when "11101110001110",
                             3279 when "11101110001111",
                             3279 when "11101110010000",
                             3279 when "11101110010001",
                             3279 when "11101110010010",
                             3278 when "11101110010011",
                             3278 when "11101110010100",
                             3278 when "11101110010101",
                             3278 when "11101110010110",
                             3278 when "11101110010111",
                             3277 when "11101110011000",
                             3277 when "11101110011001",
                             3277 when "11101110011010",
                             3277 when "11101110011011",
                             3277 when "11101110011100",
                             3276 when "11101110011101",
                             3276 when "11101110011110",
                             3276 when "11101110011111",
                             3276 when "11101110100000",
                             3275 when "11101110100001",
                             3275 when "11101110100010",
                             3275 when "11101110100011",
                             3275 when "11101110100100",
                             3275 when "11101110100101",
                             3274 when "11101110100110",
                             3274 when "11101110100111",
                             3274 when "11101110101000",
                             3274 when "11101110101001",
                             3274 when "11101110101010",
                             3273 when "11101110101011",
                             3273 when "11101110101100",
                             3273 when "11101110101101",
                             3273 when "11101110101110",
                             3272 when "11101110101111",
                             3272 when "11101110110000",
                             3272 when "11101110110001",
                             3272 when "11101110110010",
                             3272 when "11101110110011",
                             3271 when "11101110110100",
                             3271 when "11101110110101",
                             3271 when "11101110110110",
                             3271 when "11101110110111",
                             3271 when "11101110111000",
                             3270 when "11101110111001",
                             3270 when "11101110111010",
                             3270 when "11101110111011",
                             3270 when "11101110111100",
                             3269 when "11101110111101",
                             3269 when "11101110111110",
                             3269 when "11101110111111",
                             3269 when "11101111000000",
                             3269 when "11101111000001",
                             3268 when "11101111000010",
                             3268 when "11101111000011",
                             3268 when "11101111000100",
                             3268 when "11101111000101",
                             3268 when "11101111000110",
                             3267 when "11101111000111",
                             3267 when "11101111001000",
                             3267 when "11101111001001",
                             3267 when "11101111001010",
                             3266 when "11101111001011",
                             3266 when "11101111001100",
                             3266 when "11101111001101",
                             3266 when "11101111001110",
                             3266 when "11101111001111",
                             3265 when "11101111010000",
                             3265 when "11101111010001",
                             3265 when "11101111010010",
                             3265 when "11101111010011",
                             3265 when "11101111010100",
                             3264 when "11101111010101",
                             3264 when "11101111010110",
                             3264 when "11101111010111",
                             3264 when "11101111011000",
                             3263 when "11101111011001",
                             3263 when "11101111011010",
                             3263 when "11101111011011",
                             3263 when "11101111011100",
                             3263 when "11101111011101",
                             3262 when "11101111011110",
                             3262 when "11101111011111",
                             3262 when "11101111100000",
                             3262 when "11101111100001",
                             3262 when "11101111100010",
                             3261 when "11101111100011",
                             3261 when "11101111100100",
                             3261 when "11101111100101",
                             3261 when "11101111100110",
                             3261 when "11101111100111",
                             3260 when "11101111101000",
                             3260 when "11101111101001",
                             3260 when "11101111101010",
                             3260 when "11101111101011",
                             3259 when "11101111101100",
                             3259 when "11101111101101",
                             3259 when "11101111101110",
                             3259 when "11101111101111",
                             3259 when "11101111110000",
                             3258 when "11101111110001",
                             3258 when "11101111110010",
                             3258 when "11101111110011",
                             3258 when "11101111110100",
                             3258 when "11101111110101",
                             3257 when "11101111110110",
                             3257 when "11101111110111",
                             3257 when "11101111111000",
                             3257 when "11101111111001",
                             3256 when "11101111111010",
                             3256 when "11101111111011",
                             3256 when "11101111111100",
                             3256 when "11101111111101",
                             3256 when "11101111111110",
                             3255 when "11101111111111",
                             3255 when "11110000000000",
                             3255 when "11110000000001",
                             3255 when "11110000000010",
                             3255 when "11110000000011",
                             3254 when "11110000000100",
                             3254 when "11110000000101",
                             3254 when "11110000000110",
                             3254 when "11110000000111",
                             3254 when "11110000001000",
                             3253 when "11110000001001",
                             3253 when "11110000001010",
                             3253 when "11110000001011",
                             3253 when "11110000001100",
                             3252 when "11110000001101",
                             3252 when "11110000001110",
                             3252 when "11110000001111",
                             3252 when "11110000010000",
                             3252 when "11110000010001",
                             3251 when "11110000010010",
                             3251 when "11110000010011",
                             3251 when "11110000010100",
                             3251 when "11110000010101",
                             3251 when "11110000010110",
                             3250 when "11110000010111",
                             3250 when "11110000011000",
                             3250 when "11110000011001",
                             3250 when "11110000011010",
                             3249 when "11110000011011",
                             3249 when "11110000011100",
                             3249 when "11110000011101",
                             3249 when "11110000011110",
                             3249 when "11110000011111",
                             3248 when "11110000100000",
                             3248 when "11110000100001",
                             3248 when "11110000100010",
                             3248 when "11110000100011",
                             3248 when "11110000100100",
                             3247 when "11110000100101",
                             3247 when "11110000100110",
                             3247 when "11110000100111",
                             3247 when "11110000101000",
                             3247 when "11110000101001",
                             3246 when "11110000101010",
                             3246 when "11110000101011",
                             3246 when "11110000101100",
                             3246 when "11110000101101",
                             3245 when "11110000101110",
                             3245 when "11110000101111",
                             3245 when "11110000110000",
                             3245 when "11110000110001",
                             3245 when "11110000110010",
                             3244 when "11110000110011",
                             3244 when "11110000110100",
                             3244 when "11110000110101",
                             3244 when "11110000110110",
                             3244 when "11110000110111",
                             3243 when "11110000111000",
                             3243 when "11110000111001",
                             3243 when "11110000111010",
                             3243 when "11110000111011",
                             3243 when "11110000111100",
                             3242 when "11110000111101",
                             3242 when "11110000111110",
                             3242 when "11110000111111",
                             3242 when "11110001000000",
                             3241 when "11110001000001",
                             3241 when "11110001000010",
                             3241 when "11110001000011",
                             3241 when "11110001000100",
                             3241 when "11110001000101",
                             3240 when "11110001000110",
                             3240 when "11110001000111",
                             3240 when "11110001001000",
                             3240 when "11110001001001",
                             3240 when "11110001001010",
                             3239 when "11110001001011",
                             3239 when "11110001001100",
                             3239 when "11110001001101",
                             3239 when "11110001001110",
                             3239 when "11110001001111",
                             3238 when "11110001010000",
                             3238 when "11110001010001",
                             3238 when "11110001010010",
                             3238 when "11110001010011",
                             3238 when "11110001010100",
                             3237 when "11110001010101",
                             3237 when "11110001010110",
                             3237 when "11110001010111",
                             3237 when "11110001011000",
                             3236 when "11110001011001",
                             3236 when "11110001011010",
                             3236 when "11110001011011",
                             3236 when "11110001011100",
                             3236 when "11110001011101",
                             3235 when "11110001011110",
                             3235 when "11110001011111",
                             3235 when "11110001100000",
                             3235 when "11110001100001",
                             3235 when "11110001100010",
                             3234 when "11110001100011",
                             3234 when "11110001100100",
                             3234 when "11110001100101",
                             3234 when "11110001100110",
                             3234 when "11110001100111",
                             3233 when "11110001101000",
                             3233 when "11110001101001",
                             3233 when "11110001101010",
                             3233 when "11110001101011",
                             3232 when "11110001101100",
                             3232 when "11110001101101",
                             3232 when "11110001101110",
                             3232 when "11110001101111",
                             3232 when "11110001110000",
                             3231 when "11110001110001",
                             3231 when "11110001110010",
                             3231 when "11110001110011",
                             3231 when "11110001110100",
                             3231 when "11110001110101",
                             3230 when "11110001110110",
                             3230 when "11110001110111",
                             3230 when "11110001111000",
                             3230 when "11110001111001",
                             3230 when "11110001111010",
                             3229 when "11110001111011",
                             3229 when "11110001111100",
                             3229 when "11110001111101",
                             3229 when "11110001111110",
                             3229 when "11110001111111",
                             3228 when "11110010000000",
                             3228 when "11110010000001",
                             3228 when "11110010000010",
                             3228 when "11110010000011",
                             3227 when "11110010000100",
                             3227 when "11110010000101",
                             3227 when "11110010000110",
                             3227 when "11110010000111",
                             3227 when "11110010001000",
                             3226 when "11110010001001",
                             3226 when "11110010001010",
                             3226 when "11110010001011",
                             3226 when "11110010001100",
                             3226 when "11110010001101",
                             3225 when "11110010001110",
                             3225 when "11110010001111",
                             3225 when "11110010010000",
                             3225 when "11110010010001",
                             3225 when "11110010010010",
                             3224 when "11110010010011",
                             3224 when "11110010010100",
                             3224 when "11110010010101",
                             3224 when "11110010010110",
                             3224 when "11110010010111",
                             3223 when "11110010011000",
                             3223 when "11110010011001",
                             3223 when "11110010011010",
                             3223 when "11110010011011",
                             3222 when "11110010011100",
                             3222 when "11110010011101",
                             3222 when "11110010011110",
                             3222 when "11110010011111",
                             3222 when "11110010100000",
                             3221 when "11110010100001",
                             3221 when "11110010100010",
                             3221 when "11110010100011",
                             3221 when "11110010100100",
                             3221 when "11110010100101",
                             3220 when "11110010100110",
                             3220 when "11110010100111",
                             3220 when "11110010101000",
                             3220 when "11110010101001",
                             3220 when "11110010101010",
                             3219 when "11110010101011",
                             3219 when "11110010101100",
                             3219 when "11110010101101",
                             3219 when "11110010101110",
                             3219 when "11110010101111",
                             3218 when "11110010110000",
                             3218 when "11110010110001",
                             3218 when "11110010110010",
                             3218 when "11110010110011",
                             3218 when "11110010110100",
                             3217 when "11110010110101",
                             3217 when "11110010110110",
                             3217 when "11110010110111",
                             3217 when "11110010111000",
                             3216 when "11110010111001",
                             3216 when "11110010111010",
                             3216 when "11110010111011",
                             3216 when "11110010111100",
                             3216 when "11110010111101",
                             3215 when "11110010111110",
                             3215 when "11110010111111",
                             3215 when "11110011000000",
                             3215 when "11110011000001",
                             3215 when "11110011000010",
                             3214 when "11110011000011",
                             3214 when "11110011000100",
                             3214 when "11110011000101",
                             3214 when "11110011000110",
                             3214 when "11110011000111",
                             3213 when "11110011001000",
                             3213 when "11110011001001",
                             3213 when "11110011001010",
                             3213 when "11110011001011",
                             3213 when "11110011001100",
                             3212 when "11110011001101",
                             3212 when "11110011001110",
                             3212 when "11110011001111",
                             3212 when "11110011010000",
                             3212 when "11110011010001",
                             3211 when "11110011010010",
                             3211 when "11110011010011",
                             3211 when "11110011010100",
                             3211 when "11110011010101",
                             3210 when "11110011010110",
                             3210 when "11110011010111",
                             3210 when "11110011011000",
                             3210 when "11110011011001",
                             3210 when "11110011011010",
                             3209 when "11110011011011",
                             3209 when "11110011011100",
                             3209 when "11110011011101",
                             3209 when "11110011011110",
                             3209 when "11110011011111",
                             3208 when "11110011100000",
                             3208 when "11110011100001",
                             3208 when "11110011100010",
                             3208 when "11110011100011",
                             3208 when "11110011100100",
                             3207 when "11110011100101",
                             3207 when "11110011100110",
                             3207 when "11110011100111",
                             3207 when "11110011101000",
                             3207 when "11110011101001",
                             3206 when "11110011101010",
                             3206 when "11110011101011",
                             3206 when "11110011101100",
                             3206 when "11110011101101",
                             3206 when "11110011101110",
                             3205 when "11110011101111",
                             3205 when "11110011110000",
                             3205 when "11110011110001",
                             3205 when "11110011110010",
                             3205 when "11110011110011",
                             3204 when "11110011110100",
                             3204 when "11110011110101",
                             3204 when "11110011110110",
                             3204 when "11110011110111",
                             3203 when "11110011111000",
                             3203 when "11110011111001",
                             3203 when "11110011111010",
                             3203 when "11110011111011",
                             3203 when "11110011111100",
                             3202 when "11110011111101",
                             3202 when "11110011111110",
                             3202 when "11110011111111",
                             3202 when "11110100000000",
                             3202 when "11110100000001",
                             3201 when "11110100000010",
                             3201 when "11110100000011",
                             3201 when "11110100000100",
                             3201 when "11110100000101",
                             3201 when "11110100000110",
                             3200 when "11110100000111",
                             3200 when "11110100001000",
                             3200 when "11110100001001",
                             3200 when "11110100001010",
                             3200 when "11110100001011",
                             3199 when "11110100001100",
                             3199 when "11110100001101",
                             3199 when "11110100001110",
                             3199 when "11110100001111",
                             3199 when "11110100010000",
                             3198 when "11110100010001",
                             3198 when "11110100010010",
                             3198 when "11110100010011",
                             3198 when "11110100010100",
                             3198 when "11110100010101",
                             3197 when "11110100010110",
                             3197 when "11110100010111",
                             3197 when "11110100011000",
                             3197 when "11110100011001",
                             3197 when "11110100011010",
                             3196 when "11110100011011",
                             3196 when "11110100011100",
                             3196 when "11110100011101",
                             3196 when "11110100011110",
                             3196 when "11110100011111",
                             3195 when "11110100100000",
                             3195 when "11110100100001",
                             3195 when "11110100100010",
                             3195 when "11110100100011",
                             3194 when "11110100100100",
                             3194 when "11110100100101",
                             3194 when "11110100100110",
                             3194 when "11110100100111",
                             3194 when "11110100101000",
                             3193 when "11110100101001",
                             3193 when "11110100101010",
                             3193 when "11110100101011",
                             3193 when "11110100101100",
                             3193 when "11110100101101",
                             3192 when "11110100101110",
                             3192 when "11110100101111",
                             3192 when "11110100110000",
                             3192 when "11110100110001",
                             3192 when "11110100110010",
                             3191 when "11110100110011",
                             3191 when "11110100110100",
                             3191 when "11110100110101",
                             3191 when "11110100110110",
                             3191 when "11110100110111",
                             3190 when "11110100111000",
                             3190 when "11110100111001",
                             3190 when "11110100111010",
                             3190 when "11110100111011",
                             3190 when "11110100111100",
                             3189 when "11110100111101",
                             3189 when "11110100111110",
                             3189 when "11110100111111",
                             3189 when "11110101000000",
                             3189 when "11110101000001",
                             3188 when "11110101000010",
                             3188 when "11110101000011",
                             3188 when "11110101000100",
                             3188 when "11110101000101",
                             3188 when "11110101000110",
                             3187 when "11110101000111",
                             3187 when "11110101001000",
                             3187 when "11110101001001",
                             3187 when "11110101001010",
                             3187 when "11110101001011",
                             3186 when "11110101001100",
                             3186 when "11110101001101",
                             3186 when "11110101001110",
                             3186 when "11110101001111",
                             3186 when "11110101010000",
                             3185 when "11110101010001",
                             3185 when "11110101010010",
                             3185 when "11110101010011",
                             3185 when "11110101010100",
                             3185 when "11110101010101",
                             3184 when "11110101010110",
                             3184 when "11110101010111",
                             3184 when "11110101011000",
                             3184 when "11110101011001",
                             3183 when "11110101011010",
                             3183 when "11110101011011",
                             3183 when "11110101011100",
                             3183 when "11110101011101",
                             3183 when "11110101011110",
                             3182 when "11110101011111",
                             3182 when "11110101100000",
                             3182 when "11110101100001",
                             3182 when "11110101100010",
                             3182 when "11110101100011",
                             3181 when "11110101100100",
                             3181 when "11110101100101",
                             3181 when "11110101100110",
                             3181 when "11110101100111",
                             3181 when "11110101101000",
                             3180 when "11110101101001",
                             3180 when "11110101101010",
                             3180 when "11110101101011",
                             3180 when "11110101101100",
                             3180 when "11110101101101",
                             3179 when "11110101101110",
                             3179 when "11110101101111",
                             3179 when "11110101110000",
                             3179 when "11110101110001",
                             3179 when "11110101110010",
                             3178 when "11110101110011",
                             3178 when "11110101110100",
                             3178 when "11110101110101",
                             3178 when "11110101110110",
                             3178 when "11110101110111",
                             3177 when "11110101111000",
                             3177 when "11110101111001",
                             3177 when "11110101111010",
                             3177 when "11110101111011",
                             3177 when "11110101111100",
                             3176 when "11110101111101",
                             3176 when "11110101111110",
                             3176 when "11110101111111",
                             3176 when "11110110000000",
                             3176 when "11110110000001",
                             3175 when "11110110000010",
                             3175 when "11110110000011",
                             3175 when "11110110000100",
                             3175 when "11110110000101",
                             3175 when "11110110000110",
                             3174 when "11110110000111",
                             3174 when "11110110001000",
                             3174 when "11110110001001",
                             3174 when "11110110001010",
                             3174 when "11110110001011",
                             3173 when "11110110001100",
                             3173 when "11110110001101",
                             3173 when "11110110001110",
                             3173 when "11110110001111",
                             3173 when "11110110010000",
                             3172 when "11110110010001",
                             3172 when "11110110010010",
                             3172 when "11110110010011",
                             3172 when "11110110010100",
                             3172 when "11110110010101",
                             3171 when "11110110010110",
                             3171 when "11110110010111",
                             3171 when "11110110011000",
                             3171 when "11110110011001",
                             3171 when "11110110011010",
                             3170 when "11110110011011",
                             3170 when "11110110011100",
                             3170 when "11110110011101",
                             3170 when "11110110011110",
                             3170 when "11110110011111",
                             3169 when "11110110100000",
                             3169 when "11110110100001",
                             3169 when "11110110100010",
                             3169 when "11110110100011",
                             3169 when "11110110100100",
                             3168 when "11110110100101",
                             3168 when "11110110100110",
                             3168 when "11110110100111",
                             3168 when "11110110101000",
                             3168 when "11110110101001",
                             3167 when "11110110101010",
                             3167 when "11110110101011",
                             3167 when "11110110101100",
                             3167 when "11110110101101",
                             3167 when "11110110101110",
                             3166 when "11110110101111",
                             3166 when "11110110110000",
                             3166 when "11110110110001",
                             3166 when "11110110110010",
                             3166 when "11110110110011",
                             3165 when "11110110110100",
                             3165 when "11110110110101",
                             3165 when "11110110110110",
                             3165 when "11110110110111",
                             3165 when "11110110111000",
                             3164 when "11110110111001",
                             3164 when "11110110111010",
                             3164 when "11110110111011",
                             3164 when "11110110111100",
                             3164 when "11110110111101",
                             3163 when "11110110111110",
                             3163 when "11110110111111",
                             3163 when "11110111000000",
                             3163 when "11110111000001",
                             3163 when "11110111000010",
                             3162 when "11110111000011",
                             3162 when "11110111000100",
                             3162 when "11110111000101",
                             3162 when "11110111000110",
                             3162 when "11110111000111",
                             3161 when "11110111001000",
                             3161 when "11110111001001",
                             3161 when "11110111001010",
                             3161 when "11110111001011",
                             3161 when "11110111001100",
                             3160 when "11110111001101",
                             3160 when "11110111001110",
                             3160 when "11110111001111",
                             3160 when "11110111010000",
                             3160 when "11110111010001",
                             3159 when "11110111010010",
                             3159 when "11110111010011",
                             3159 when "11110111010100",
                             3159 when "11110111010101",
                             3159 when "11110111010110",
                             3158 when "11110111010111",
                             3158 when "11110111011000",
                             3158 when "11110111011001",
                             3158 when "11110111011010",
                             3158 when "11110111011011",
                             3157 when "11110111011100",
                             3157 when "11110111011101",
                             3157 when "11110111011110",
                             3157 when "11110111011111",
                             3157 when "11110111100000",
                             3156 when "11110111100001",
                             3156 when "11110111100010",
                             3156 when "11110111100011",
                             3156 when "11110111100100",
                             3156 when "11110111100101",
                             3155 when "11110111100110",
                             3155 when "11110111100111",
                             3155 when "11110111101000",
                             3155 when "11110111101001",
                             3155 when "11110111101010",
                             3154 when "11110111101011",
                             3154 when "11110111101100",
                             3154 when "11110111101101",
                             3154 when "11110111101110",
                             3154 when "11110111101111",
                             3153 when "11110111110000",
                             3153 when "11110111110001",
                             3153 when "11110111110010",
                             3153 when "11110111110011",
                             3153 when "11110111110100",
                             3152 when "11110111110101",
                             3152 when "11110111110110",
                             3152 when "11110111110111",
                             3152 when "11110111111000",
                             3152 when "11110111111001",
                             3151 when "11110111111010",
                             3151 when "11110111111011",
                             3151 when "11110111111100",
                             3151 when "11110111111101",
                             3151 when "11110111111110",
                             3150 when "11110111111111",
                             3150 when "11111000000000",
                             3150 when "11111000000001",
                             3150 when "11111000000010",
                             3150 when "11111000000011",
                             3149 when "11111000000100",
                             3149 when "11111000000101",
                             3149 when "11111000000110",
                             3149 when "11111000000111",
                             3149 when "11111000001000",
                             3148 when "11111000001001",
                             3148 when "11111000001010",
                             3148 when "11111000001011",
                             3148 when "11111000001100",
                             3148 when "11111000001101",
                             3147 when "11111000001110",
                             3147 when "11111000001111",
                             3147 when "11111000010000",
                             3147 when "11111000010001",
                             3147 when "11111000010010",
                             3146 when "11111000010011",
                             3146 when "11111000010100",
                             3146 when "11111000010101",
                             3146 when "11111000010110",
                             3146 when "11111000010111",
                             3145 when "11111000011000",
                             3145 when "11111000011001",
                             3145 when "11111000011010",
                             3145 when "11111000011011",
                             3145 when "11111000011100",
                             3144 when "11111000011101",
                             3144 when "11111000011110",
                             3144 when "11111000011111",
                             3144 when "11111000100000",
                             3144 when "11111000100001",
                             3143 when "11111000100010",
                             3143 when "11111000100011",
                             3143 when "11111000100100",
                             3143 when "11111000100101",
                             3143 when "11111000100110",
                             3142 when "11111000100111",
                             3142 when "11111000101000",
                             3142 when "11111000101001",
                             3142 when "11111000101010",
                             3142 when "11111000101011",
                             3141 when "11111000101100",
                             3141 when "11111000101101",
                             3141 when "11111000101110",
                             3141 when "11111000101111",
                             3141 when "11111000110000",
                             3141 when "11111000110001",
                             3140 when "11111000110010",
                             3140 when "11111000110011",
                             3140 when "11111000110100",
                             3140 when "11111000110101",
                             3140 when "11111000110110",
                             3139 when "11111000110111",
                             3139 when "11111000111000",
                             3139 when "11111000111001",
                             3139 when "11111000111010",
                             3139 when "11111000111011",
                             3138 when "11111000111100",
                             3138 when "11111000111101",
                             3138 when "11111000111110",
                             3138 when "11111000111111",
                             3138 when "11111001000000",
                             3137 when "11111001000001",
                             3137 when "11111001000010",
                             3137 when "11111001000011",
                             3137 when "11111001000100",
                             3137 when "11111001000101",
                             3136 when "11111001000110",
                             3136 when "11111001000111",
                             3136 when "11111001001000",
                             3136 when "11111001001001",
                             3136 when "11111001001010",
                             3135 when "11111001001011",
                             3135 when "11111001001100",
                             3135 when "11111001001101",
                             3135 when "11111001001110",
                             3135 when "11111001001111",
                             3134 when "11111001010000",
                             3134 when "11111001010001",
                             3134 when "11111001010010",
                             3134 when "11111001010011",
                             3134 when "11111001010100",
                             3133 when "11111001010101",
                             3133 when "11111001010110",
                             3133 when "11111001010111",
                             3133 when "11111001011000",
                             3133 when "11111001011001",
                             3132 when "11111001011010",
                             3132 when "11111001011011",
                             3132 when "11111001011100",
                             3132 when "11111001011101",
                             3132 when "11111001011110",
                             3131 when "11111001011111",
                             3131 when "11111001100000",
                             3131 when "11111001100001",
                             3131 when "11111001100010",
                             3131 when "11111001100011",
                             3130 when "11111001100100",
                             3130 when "11111001100101",
                             3130 when "11111001100110",
                             3130 when "11111001100111",
                             3130 when "11111001101000",
                             3129 when "11111001101001",
                             3129 when "11111001101010",
                             3129 when "11111001101011",
                             3129 when "11111001101100",
                             3129 when "11111001101101",
                             3129 when "11111001101110",
                             3128 when "11111001101111",
                             3128 when "11111001110000",
                             3128 when "11111001110001",
                             3128 when "11111001110010",
                             3128 when "11111001110011",
                             3127 when "11111001110100",
                             3127 when "11111001110101",
                             3127 when "11111001110110",
                             3127 when "11111001110111",
                             3127 when "11111001111000",
                             3126 when "11111001111001",
                             3126 when "11111001111010",
                             3126 when "11111001111011",
                             3126 when "11111001111100",
                             3126 when "11111001111101",
                             3125 when "11111001111110",
                             3125 when "11111001111111",
                             3125 when "11111010000000",
                             3125 when "11111010000001",
                             3125 when "11111010000010",
                             3124 when "11111010000011",
                             3124 when "11111010000100",
                             3124 when "11111010000101",
                             3124 when "11111010000110",
                             3124 when "11111010000111",
                             3123 when "11111010001000",
                             3123 when "11111010001001",
                             3123 when "11111010001010",
                             3123 when "11111010001011",
                             3123 when "11111010001100",
                             3122 when "11111010001101",
                             3122 when "11111010001110",
                             3122 when "11111010001111",
                             3122 when "11111010010000",
                             3122 when "11111010010001",
                             3121 when "11111010010010",
                             3121 when "11111010010011",
                             3121 when "11111010010100",
                             3121 when "11111010010101",
                             3121 when "11111010010110",
                             3121 when "11111010010111",
                             3120 when "11111010011000",
                             3120 when "11111010011001",
                             3120 when "11111010011010",
                             3120 when "11111010011011",
                             3120 when "11111010011100",
                             3119 when "11111010011101",
                             3119 when "11111010011110",
                             3119 when "11111010011111",
                             3119 when "11111010100000",
                             3119 when "11111010100001",
                             3118 when "11111010100010",
                             3118 when "11111010100011",
                             3118 when "11111010100100",
                             3118 when "11111010100101",
                             3118 when "11111010100110",
                             3117 when "11111010100111",
                             3117 when "11111010101000",
                             3117 when "11111010101001",
                             3117 when "11111010101010",
                             3117 when "11111010101011",
                             3116 when "11111010101100",
                             3116 when "11111010101101",
                             3116 when "11111010101110",
                             3116 when "11111010101111",
                             3116 when "11111010110000",
                             3115 when "11111010110001",
                             3115 when "11111010110010",
                             3115 when "11111010110011",
                             3115 when "11111010110100",
                             3115 when "11111010110101",
                             3114 when "11111010110110",
                             3114 when "11111010110111",
                             3114 when "11111010111000",
                             3114 when "11111010111001",
                             3114 when "11111010111010",
                             3114 when "11111010111011",
                             3113 when "11111010111100",
                             3113 when "11111010111101",
                             3113 when "11111010111110",
                             3113 when "11111010111111",
                             3113 when "11111011000000",
                             3112 when "11111011000001",
                             3112 when "11111011000010",
                             3112 when "11111011000011",
                             3112 when "11111011000100",
                             3112 when "11111011000101",
                             3111 when "11111011000110",
                             3111 when "11111011000111",
                             3111 when "11111011001000",
                             3111 when "11111011001001",
                             3111 when "11111011001010",
                             3110 when "11111011001011",
                             3110 when "11111011001100",
                             3110 when "11111011001101",
                             3110 when "11111011001110",
                             3110 when "11111011001111",
                             3109 when "11111011010000",
                             3109 when "11111011010001",
                             3109 when "11111011010010",
                             3109 when "11111011010011",
                             3109 when "11111011010100",
                             3108 when "11111011010101",
                             3108 when "11111011010110",
                             3108 when "11111011010111",
                             3108 when "11111011011000",
                             3108 when "11111011011001",
                             3108 when "11111011011010",
                             3107 when "11111011011011",
                             3107 when "11111011011100",
                             3107 when "11111011011101",
                             3107 when "11111011011110",
                             3107 when "11111011011111",
                             3106 when "11111011100000",
                             3106 when "11111011100001",
                             3106 when "11111011100010",
                             3106 when "11111011100011",
                             3106 when "11111011100100",
                             3105 when "11111011100101",
                             3105 when "11111011100110",
                             3105 when "11111011100111",
                             3105 when "11111011101000",
                             3105 when "11111011101001",
                             3104 when "11111011101010",
                             3104 when "11111011101011",
                             3104 when "11111011101100",
                             3104 when "11111011101101",
                             3104 when "11111011101110",
                             3103 when "11111011101111",
                             3103 when "11111011110000",
                             3103 when "11111011110001",
                             3103 when "11111011110010",
                             3103 when "11111011110011",
                             3103 when "11111011110100",
                             3102 when "11111011110101",
                             3102 when "11111011110110",
                             3102 when "11111011110111",
                             3102 when "11111011111000",
                             3102 when "11111011111001",
                             3101 when "11111011111010",
                             3101 when "11111011111011",
                             3101 when "11111011111100",
                             3101 when "11111011111101",
                             3101 when "11111011111110",
                             3100 when "11111011111111",
                             3100 when "11111100000000",
                             3100 when "11111100000001",
                             3100 when "11111100000010",
                             3100 when "11111100000011",
                             3099 when "11111100000100",
                             3099 when "11111100000101",
                             3099 when "11111100000110",
                             3099 when "11111100000111",
                             3099 when "11111100001000",
                             3098 when "11111100001001",
                             3098 when "11111100001010",
                             3098 when "11111100001011",
                             3098 when "11111100001100",
                             3098 when "11111100001101",
                             3098 when "11111100001110",
                             3097 when "11111100001111",
                             3097 when "11111100010000",
                             3097 when "11111100010001",
                             3097 when "11111100010010",
                             3097 when "11111100010011",
                             3096 when "11111100010100",
                             3096 when "11111100010101",
                             3096 when "11111100010110",
                             3096 when "11111100010111",
                             3096 when "11111100011000",
                             3095 when "11111100011001",
                             3095 when "11111100011010",
                             3095 when "11111100011011",
                             3095 when "11111100011100",
                             3095 when "11111100011101",
                             3094 when "11111100011110",
                             3094 when "11111100011111",
                             3094 when "11111100100000",
                             3094 when "11111100100001",
                             3094 when "11111100100010",
                             3093 when "11111100100011",
                             3093 when "11111100100100",
                             3093 when "11111100100101",
                             3093 when "11111100100110",
                             3093 when "11111100100111",
                             3093 when "11111100101000",
                             3092 when "11111100101001",
                             3092 when "11111100101010",
                             3092 when "11111100101011",
                             3092 when "11111100101100",
                             3092 when "11111100101101",
                             3091 when "11111100101110",
                             3091 when "11111100101111",
                             3091 when "11111100110000",
                             3091 when "11111100110001",
                             3091 when "11111100110010",
                             3090 when "11111100110011",
                             3090 when "11111100110100",
                             3090 when "11111100110101",
                             3090 when "11111100110110",
                             3090 when "11111100110111",
                             3089 when "11111100111000",
                             3089 when "11111100111001",
                             3089 when "11111100111010",
                             3089 when "11111100111011",
                             3089 when "11111100111100",
                             3089 when "11111100111101",
                             3088 when "11111100111110",
                             3088 when "11111100111111",
                             3088 when "11111101000000",
                             3088 when "11111101000001",
                             3088 when "11111101000010",
                             3087 when "11111101000011",
                             3087 when "11111101000100",
                             3087 when "11111101000101",
                             3087 when "11111101000110",
                             3087 when "11111101000111",
                             3086 when "11111101001000",
                             3086 when "11111101001001",
                             3086 when "11111101001010",
                             3086 when "11111101001011",
                             3086 when "11111101001100",
                             3085 when "11111101001101",
                             3085 when "11111101001110",
                             3085 when "11111101001111",
                             3085 when "11111101010000",
                             3085 when "11111101010001",
                             3085 when "11111101010010",
                             3084 when "11111101010011",
                             3084 when "11111101010100",
                             3084 when "11111101010101",
                             3084 when "11111101010110",
                             3084 when "11111101010111",
                             3083 when "11111101011000",
                             3083 when "11111101011001",
                             3083 when "11111101011010",
                             3083 when "11111101011011",
                             3083 when "11111101011100",
                             3082 when "11111101011101",
                             3082 when "11111101011110",
                             3082 when "11111101011111",
                             3082 when "11111101100000",
                             3082 when "11111101100001",
                             3081 when "11111101100010",
                             3081 when "11111101100011",
                             3081 when "11111101100100",
                             3081 when "11111101100101",
                             3081 when "11111101100110",
                             3081 when "11111101100111",
                             3080 when "11111101101000",
                             3080 when "11111101101001",
                             3080 when "11111101101010",
                             3080 when "11111101101011",
                             3080 when "11111101101100",
                             3079 when "11111101101101",
                             3079 when "11111101101110",
                             3079 when "11111101101111",
                             3079 when "11111101110000",
                             3079 when "11111101110001",
                             3078 when "11111101110010",
                             3078 when "11111101110011",
                             3078 when "11111101110100",
                             3078 when "11111101110101",
                             3078 when "11111101110110",
                             3077 when "11111101110111",
                             3077 when "11111101111000",
                             3077 when "11111101111001",
                             3077 when "11111101111010",
                             3077 when "11111101111011",
                             3077 when "11111101111100",
                             3076 when "11111101111101",
                             3076 when "11111101111110",
                             3076 when "11111101111111",
                             3076 when "11111110000000",
                             3076 when "11111110000001",
                             3075 when "11111110000010",
                             3075 when "11111110000011",
                             3075 when "11111110000100",
                             3075 when "11111110000101",
                             3075 when "11111110000110",
                             3074 when "11111110000111",
                             3074 when "11111110001000",
                             3074 when "11111110001001",
                             3074 when "11111110001010",
                             3074 when "11111110001011",
                             3074 when "11111110001100",
                             3073 when "11111110001101",
                             3073 when "11111110001110",
                             3073 when "11111110001111",
                             3073 when "11111110010000",
                             3073 when "11111110010001",
                             3072 when "11111110010010",
                             3072 when "11111110010011",
                             3072 when "11111110010100",
                             3072 when "11111110010101",
                             3072 when "11111110010110",
                             3071 when "11111110010111",
                             3071 when "11111110011000",
                             3071 when "11111110011001",
                             3071 when "11111110011010",
                             3071 when "11111110011011",
                             3070 when "11111110011100",
                             3070 when "11111110011101",
                             3070 when "11111110011110",
                             3070 when "11111110011111",
                             3070 when "11111110100000",
                             3070 when "11111110100001",
                             3069 when "11111110100010",
                             3069 when "11111110100011",
                             3069 when "11111110100100",
                             3069 when "11111110100101",
                             3069 when "11111110100110",
                             3068 when "11111110100111",
                             3068 when "11111110101000",
                             3068 when "11111110101001",
                             3068 when "11111110101010",
                             3068 when "11111110101011",
                             3067 when "11111110101100",
                             3067 when "11111110101101",
                             3067 when "11111110101110",
                             3067 when "11111110101111",
                             3067 when "11111110110000",
                             3067 when "11111110110001",
                             3066 when "11111110110010",
                             3066 when "11111110110011",
                             3066 when "11111110110100",
                             3066 when "11111110110101",
                             3066 when "11111110110110",
                             3065 when "11111110110111",
                             3065 when "11111110111000",
                             3065 when "11111110111001",
                             3065 when "11111110111010",
                             3065 when "11111110111011",
                             3064 when "11111110111100",
                             3064 when "11111110111101",
                             3064 when "11111110111110",
                             3064 when "11111110111111",
                             3064 when "11111111000000",
                             3064 when "11111111000001",
                             3063 when "11111111000010",
                             3063 when "11111111000011",
                             3063 when "11111111000100",
                             3063 when "11111111000101",
                             3063 when "11111111000110",
                             3062 when "11111111000111",
                             3062 when "11111111001000",
                             3062 when "11111111001001",
                             3062 when "11111111001010",
                             3062 when "11111111001011",
                             3061 when "11111111001100",
                             3061 when "11111111001101",
                             3061 when "11111111001110",
                             3061 when "11111111001111",
                             3061 when "11111111010000",
                             3061 when "11111111010001",
                             3060 when "11111111010010",
                             3060 when "11111111010011",
                             3060 when "11111111010100",
                             3060 when "11111111010101",
                             3060 when "11111111010110",
                             3059 when "11111111010111",
                             3059 when "11111111011000",
                             3059 when "11111111011001",
                             3059 when "11111111011010",
                             3059 when "11111111011011",
                             3058 when "11111111011100",
                             3058 when "11111111011101",
                             3058 when "11111111011110",
                             3058 when "11111111011111",
                             3058 when "11111111100000",
                             3058 when "11111111100001",
                             3057 when "11111111100010",
                             3057 when "11111111100011",
                             3057 when "11111111100100",
                             3057 when "11111111100101",
                             3057 when "11111111100110",
                             3056 when "11111111100111",
                             3056 when "11111111101000",
                             3056 when "11111111101001",
                             3056 when "11111111101010",
                             3056 when "11111111101011",
                             3055 when "11111111101100",
                             3055 when "11111111101101",
                             3055 when "11111111101110",
                             3055 when "11111111101111",
                             3055 when "11111111110000",
                             3055 when "11111111110001",
                             3054 when "11111111110010",
                             3054 when "11111111110011",
                             3054 when "11111111110100",
                             3054 when "11111111110101",
                             3054 when "11111111110110",
                             3053 when "11111111110111",
                             3053 when "11111111111000",
                             3053 when "11111111111001",
                             3053 when "11111111111010",
                             3053 when "11111111111011",
                             3053 when "11111111111100",
                             3052 when "11111111111101",
                             3052 when "11111111111110",
                             3052 when "11111111111111",
                             0 when others;
end Behavioral;
