-- Keelin Becker-Wheeler
-- lut_sine_mem_addr.vhd

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

entity lut_sine_mem_addr is
    port (
        freq            : in  std_logic_vector(13 downto 0);
        nine_incr_ticks : out integer
    );
end lut_sine_mem_addr;

architecture Behavioral of lut_sine_mem_addr is
begin

with freq select
  nine_incr_ticks <=  0 when "00000000000000",
                      219727 when "00000000000001",
                      109863 when "00000000000010",
                      73242 when "00000000000011",
                      54932 when "00000000000100",
                      43945 when "00000000000101",
                      36621 when "00000000000110",
                      31390 when "00000000000111",
                      27466 when "00000000001000",
                      24414 when "00000000001001",
                      21973 when "00000000001010",
                      19975 when "00000000001011",
                      18311 when "00000000001100",
                      16902 when "00000000001101",
                      15695 when "00000000001110",
                      14648 when "00000000001111",
                      13733 when "00000000010000",
                      12925 when "00000000010001",
                      12207 when "00000000010010",
                      11565 when "00000000010011",
                      10986 when "00000000010100",
                      10463 when "00000000010101",
                      9988 when "00000000010110",
                      9553 when "00000000010111",
                      9155 when "00000000011000",
                      8789 when "00000000011001",
                      8451 when "00000000011010",
                      8138 when "00000000011011",
                      7847 when "00000000011100",
                      7577 when "00000000011101",
                      7324 when "00000000011110",
                      7088 when "00000000011111",
                      6866 when "00000000100000",
                      6658 when "00000000100001",
                      6463 when "00000000100010",
                      6278 when "00000000100011",
                      6104 when "00000000100100",
                      5939 when "00000000100101",
                      5782 when "00000000100110",
                      5634 when "00000000100111",
                      5493 when "00000000101000",
                      5359 when "00000000101001",
                      5232 when "00000000101010",
                      5110 when "00000000101011",
                      4994 when "00000000101100",
                      4883 when "00000000101101",
                      4777 when "00000000101110",
                      4675 when "00000000101111",
                      4578 when "00000000110000",
                      4484 when "00000000110001",
                      4395 when "00000000110010",
                      4308 when "00000000110011",
                      4226 when "00000000110100",
                      4146 when "00000000110101",
                      4069 when "00000000110110",
                      3995 when "00000000110111",
                      3924 when "00000000111000",
                      3855 when "00000000111001",
                      3788 when "00000000111010",
                      3724 when "00000000111011",
                      3662 when "00000000111100",
                      3602 when "00000000111101",
                      3544 when "00000000111110",
                      3488 when "00000000111111",
                      3433 when "00000001000000",
                      3380 when "00000001000001",
                      3329 when "00000001000010",
                      3280 when "00000001000011",
                      3231 when "00000001000100",
                      3184 when "00000001000101",
                      3139 when "00000001000110",
                      3095 when "00000001000111",
                      3052 when "00000001001000",
                      3010 when "00000001001001",
                      2969 when "00000001001010",
                      2930 when "00000001001011",
                      2891 when "00000001001100",
                      2854 when "00000001001101",
                      2817 when "00000001001110",
                      2781 when "00000001001111",
                      2747 when "00000001010000",
                      2713 when "00000001010001",
                      2680 when "00000001010010",
                      2647 when "00000001010011",
                      2616 when "00000001010100",
                      2585 when "00000001010101",
                      2555 when "00000001010110",
                      2526 when "00000001010111",
                      2497 when "00000001011000",
                      2469 when "00000001011001",
                      2441 when "00000001011010",
                      2415 when "00000001011011",
                      2388 when "00000001011100",
                      2363 when "00000001011101",
                      2338 when "00000001011110",
                      2313 when "00000001011111",
                      2289 when "00000001100000",
                      2265 when "00000001100001",
                      2242 when "00000001100010",
                      2219 when "00000001100011",
                      2197 when "00000001100100",
                      2176 when "00000001100101",
                      2154 when "00000001100110",
                      2133 when "00000001100111",
                      2113 when "00000001101000",
                      2093 when "00000001101001",
                      2073 when "00000001101010",
                      2054 when "00000001101011",
                      2035 when "00000001101100",
                      2016 when "00000001101101",
                      1998 when "00000001101110",
                      1980 when "00000001101111",
                      1962 when "00000001110000",
                      1944 when "00000001110001",
                      1927 when "00000001110010",
                      1911 when "00000001110011",
                      1894 when "00000001110100",
                      1878 when "00000001110101",
                      1862 when "00000001110110",
                      1846 when "00000001110111",
                      1831 when "00000001111000",
                      1816 when "00000001111001",
                      1801 when "00000001111010",
                      1786 when "00000001111011",
                      1772 when "00000001111100",
                      1758 when "00000001111101",
                      1744 when "00000001111110",
                      1730 when "00000001111111",
                      1717 when "00000010000000",
                      1703 when "00000010000001",
                      1690 when "00000010000010",
                      1677 when "00000010000011",
                      1665 when "00000010000100",
                      1652 when "00000010000101",
                      1640 when "00000010000110",
                      1628 when "00000010000111",
                      1616 when "00000010001000",
                      1604 when "00000010001001",
                      1592 when "00000010001010",
                      1581 when "00000010001011",
                      1569 when "00000010001100",
                      1558 when "00000010001101",
                      1547 when "00000010001110",
                      1537 when "00000010001111",
                      1526 when "00000010010000",
                      1515 when "00000010010001",
                      1505 when "00000010010010",
                      1495 when "00000010010011",
                      1485 when "00000010010100",
                      1475 when "00000010010101",
                      1465 when "00000010010110",
                      1455 when "00000010010111",
                      1446 when "00000010011000",
                      1436 when "00000010011001",
                      1427 when "00000010011010",
                      1418 when "00000010011011",
                      1409 when "00000010011100",
                      1400 when "00000010011101",
                      1391 when "00000010011110",
                      1382 when "00000010011111",
                      1373 when "00000010100000",
                      1365 when "00000010100001",
                      1356 when "00000010100010",
                      1348 when "00000010100011",
                      1340 when "00000010100100",
                      1332 when "00000010100101",
                      1324 when "00000010100110",
                      1316 when "00000010100111",
                      1308 when "00000010101000",
                      1300 when "00000010101001",
                      1293 when "00000010101010",
                      1285 when "00000010101011",
                      1277 when "00000010101100",
                      1270 when "00000010101101",
                      1263 when "00000010101110",
                      1256 when "00000010101111",
                      1248 when "00000010110000",
                      1241 when "00000010110001",
                      1234 when "00000010110010",
                      1228 when "00000010110011",
                      1221 when "00000010110100",
                      1214 when "00000010110101",
                      1207 when "00000010110110",
                      1201 when "00000010110111",
                      1194 when "00000010111000",
                      1188 when "00000010111001",
                      1181 when "00000010111010",
                      1175 when "00000010111011",
                      1169 when "00000010111100",
                      1163 when "00000010111101",
                      1156 when "00000010111110",
                      1150 when "00000010111111",
                      1144 when "00000011000000",
                      1138 when "00000011000001",
                      1133 when "00000011000010",
                      1127 when "00000011000011",
                      1121 when "00000011000100",
                      1115 when "00000011000101",
                      1110 when "00000011000110",
                      1104 when "00000011000111",
                      1099 when "00000011001000",
                      1093 when "00000011001001",
                      1088 when "00000011001010",
                      1082 when "00000011001011",
                      1077 when "00000011001100",
                      1072 when "00000011001101",
                      1067 when "00000011001110",
                      1061 when "00000011001111",
                      1056 when "00000011010000",
                      1051 when "00000011010001",
                      1046 when "00000011010010",
                      1041 when "00000011010011",
                      1036 when "00000011010100",
                      1032 when "00000011010101",
                      1027 when "00000011010110",
                      1022 when "00000011010111",
                      1017 when "00000011011000",
                      1013 when "00000011011001",
                      1008 when "00000011011010",
                      1003 when "00000011011011",
                      999 when "00000011011100",
                      994 when "00000011011101",
                      990 when "00000011011110",
                      985 when "00000011011111",
                      981 when "00000011100000",
                      977 when "00000011100001",
                      972 when "00000011100010",
                      968 when "00000011100011",
                      964 when "00000011100100",
                      960 when "00000011100101",
                      955 when "00000011100110",
                      951 when "00000011100111",
                      947 when "00000011101000",
                      943 when "00000011101001",
                      939 when "00000011101010",
                      935 when "00000011101011",
                      931 when "00000011101100",
                      927 when "00000011101101",
                      923 when "00000011101110",
                      919 when "00000011101111",
                      916 when "00000011110000",
                      912 when "00000011110001",
                      908 when "00000011110010",
                      904 when "00000011110011",
                      901 when "00000011110100",
                      897 when "00000011110101",
                      893 when "00000011110110",
                      890 when "00000011110111",
                      886 when "00000011111000",
                      882 when "00000011111001",
                      879 when "00000011111010",
                      875 when "00000011111011",
                      872 when "00000011111100",
                      868 when "00000011111101",
                      865 when "00000011111110",
                      862 when "00000011111111",
                      858 when "00000100000000",
                      855 when "00000100000001",
                      852 when "00000100000010",
                      848 when "00000100000011",
                      845 when "00000100000100",
                      842 when "00000100000101",
                      839 when "00000100000110",
                      835 when "00000100000111",
                      832 when "00000100001000",
                      829 when "00000100001001",
                      826 when "00000100001010",
                      823 when "00000100001011",
                      820 when "00000100001100",
                      817 when "00000100001101",
                      814 when "00000100001110",
                      811 when "00000100001111",
                      808 when "00000100010000",
                      805 when "00000100010001",
                      802 when "00000100010010",
                      799 when "00000100010011",
                      796 when "00000100010100",
                      793 when "00000100010101",
                      790 when "00000100010110",
                      788 when "00000100010111",
                      785 when "00000100011000",
                      782 when "00000100011001",
                      779 when "00000100011010",
                      776 when "00000100011011",
                      774 when "00000100011100",
                      771 when "00000100011101",
                      768 when "00000100011110",
                      766 when "00000100011111",
                      763 when "00000100100000",
                      760 when "00000100100001",
                      758 when "00000100100010",
                      755 when "00000100100011",
                      752 when "00000100100100",
                      750 when "00000100100101",
                      747 when "00000100100110",
                      745 when "00000100100111",
                      742 when "00000100101000",
                      740 when "00000100101001",
                      737 when "00000100101010",
                      735 when "00000100101011",
                      732 when "00000100101100",
                      730 when "00000100101101",
                      728 when "00000100101110",
                      725 when "00000100101111",
                      723 when "00000100110000",
                      720 when "00000100110001",
                      718 when "00000100110010",
                      716 when "00000100110011",
                      713 when "00000100110100",
                      711 when "00000100110101",
                      709 when "00000100110110",
                      707 when "00000100110111",
                      704 when "00000100111000",
                      702 when "00000100111001",
                      700 when "00000100111010",
                      698 when "00000100111011",
                      695 when "00000100111100",
                      693 when "00000100111101",
                      691 when "00000100111110",
                      689 when "00000100111111",
                      687 when "00000101000000",
                      685 when "00000101000001",
                      682 when "00000101000010",
                      680 when "00000101000011",
                      678 when "00000101000100",
                      676 when "00000101000101",
                      674 when "00000101000110",
                      672 when "00000101000111",
                      670 when "00000101001000",
                      668 when "00000101001001",
                      666 when "00000101001010",
                      664 when "00000101001011",
                      662 when "00000101001100",
                      660 when "00000101001101",
                      658 when "00000101001110",
                      656 when "00000101001111",
                      654 when "00000101010000",
                      652 when "00000101010001",
                      650 when "00000101010010",
                      648 when "00000101010011",
                      646 when "00000101010100",
                      644 when "00000101010101",
                      642 when "00000101010110",
                      641 when "00000101010111",
                      639 when "00000101011000",
                      637 when "00000101011001",
                      635 when "00000101011010",
                      633 when "00000101011011",
                      631 when "00000101011100",
                      630 when "00000101011101",
                      628 when "00000101011110",
                      626 when "00000101011111",
                      624 when "00000101100000",
                      622 when "00000101100001",
                      621 when "00000101100010",
                      619 when "00000101100011",
                      617 when "00000101100100",
                      615 when "00000101100101",
                      614 when "00000101100110",
                      612 when "00000101100111",
                      610 when "00000101101000",
                      609 when "00000101101001",
                      607 when "00000101101010",
                      605 when "00000101101011",
                      604 when "00000101101100",
                      602 when "00000101101101",
                      600 when "00000101101110",
                      599 when "00000101101111",
                      597 when "00000101110000",
                      595 when "00000101110001",
                      594 when "00000101110010",
                      592 when "00000101110011",
                      591 when "00000101110100",
                      589 when "00000101110101",
                      588 when "00000101110110",
                      586 when "00000101110111",
                      584 when "00000101111000",
                      583 when "00000101111001",
                      581 when "00000101111010",
                      580 when "00000101111011",
                      578 when "00000101111100",
                      577 when "00000101111101",
                      575 when "00000101111110",
                      574 when "00000101111111",
                      572 when "00000110000000",
                      571 when "00000110000001",
                      569 when "00000110000010",
                      568 when "00000110000011",
                      566 when "00000110000100",
                      565 when "00000110000101",
                      563 when "00000110000110",
                      562 when "00000110000111",
                      561 when "00000110001000",
                      559 when "00000110001001",
                      558 when "00000110001010",
                      556 when "00000110001011",
                      555 when "00000110001100",
                      553 when "00000110001101",
                      552 when "00000110001110",
                      551 when "00000110001111",
                      549 when "00000110010000",
                      548 when "00000110010001",
                      547 when "00000110010010",
                      545 when "00000110010011",
                      544 when "00000110010100",
                      543 when "00000110010101",
                      541 when "00000110010110",
                      540 when "00000110010111",
                      539 when "00000110011000",
                      537 when "00000110011001",
                      536 when "00000110011010",
                      535 when "00000110011011",
                      533 when "00000110011100",
                      532 when "00000110011101",
                      531 when "00000110011110",
                      529 when "00000110011111",
                      528 when "00000110100000",
                      527 when "00000110100001",
                      526 when "00000110100010",
                      524 when "00000110100011",
                      523 when "00000110100100",
                      522 when "00000110100101",
                      521 when "00000110100110",
                      519 when "00000110100111",
                      518 when "00000110101000",
                      517 when "00000110101001",
                      516 when "00000110101010",
                      515 when "00000110101011",
                      513 when "00000110101100",
                      512 when "00000110101101",
                      511 when "00000110101110",
                      510 when "00000110101111",
                      509 when "00000110110000",
                      507 when "00000110110001",
                      506 when "00000110110010",
                      505 when "00000110110011",
                      504 when "00000110110100",
                      503 when "00000110110101",
                      502 when "00000110110110",
                      501 when "00000110110111",
                      499 when "00000110111000",
                      498 when "00000110111001",
                      497 when "00000110111010",
                      496 when "00000110111011",
                      495 when "00000110111100",
                      494 when "00000110111101",
                      493 when "00000110111110",
                      492 when "00000110111111",
                      490 when "00000111000000",
                      489 when "00000111000001",
                      488 when "00000111000010",
                      487 when "00000111000011",
                      486 when "00000111000100",
                      485 when "00000111000101",
                      484 when "00000111000110",
                      483 when "00000111000111",
                      482 when "00000111001000",
                      481 when "00000111001001",
                      480 when "00000111001010",
                      479 when "00000111001011",
                      478 when "00000111001100",
                      477 when "00000111001101",
                      476 when "00000111001110",
                      475 when "00000111001111",
                      474 when "00000111010000",
                      473 when "00000111010001",
                      472 when "00000111010010",
                      471 when "00000111010011",
                      470 when "00000111010100",
                      469 when "00000111010101",
                      468 when "00000111010110",
                      467 when "00000111010111",
                      466 when "00000111011000",
                      465 when "00000111011001",
                      464 when "00000111011010",
                      463 when "00000111011011",
                      462 when "00000111011100",
                      461 when "00000111011101",
                      460 when "00000111011110",
                      459 when "00000111011111",
                      458 when "00000111100000",
                      457 when "00000111100001",
                      456 when "00000111100010",
                      455 when "00000111100011",
                      454 when "00000111100100",
                      453 when "00000111100101",
                      452 when "00000111100110",
                      451 when "00000111100111",
                      450 when "00000111101000",
                      449 when "00000111101001",
                      448 when "00000111101010",
                      448 when "00000111101011",
                      447 when "00000111101100",
                      446 when "00000111101101",
                      445 when "00000111101110",
                      444 when "00000111101111",
                      443 when "00000111110000",
                      442 when "00000111110001",
                      441 when "00000111110010",
                      440 when "00000111110011",
                      439 when "00000111110100",
                      439 when "00000111110101",
                      438 when "00000111110110",
                      437 when "00000111110111",
                      436 when "00000111111000",
                      435 when "00000111111001",
                      434 when "00000111111010",
                      433 when "00000111111011",
                      433 when "00000111111100",
                      432 when "00000111111101",
                      431 when "00000111111110",
                      430 when "00000111111111",
                      429 when "00001000000000",
                      428 when "00001000000001",
                      427 when "00001000000010",
                      427 when "00001000000011",
                      426 when "00001000000100",
                      425 when "00001000000101",
                      424 when "00001000000110",
                      423 when "00001000000111",
                      423 when "00001000001000",
                      422 when "00001000001001",
                      421 when "00001000001010",
                      420 when "00001000001011",
                      419 when "00001000001100",
                      419 when "00001000001101",
                      418 when "00001000001110",
                      417 when "00001000001111",
                      416 when "00001000010000",
                      415 when "00001000010001",
                      415 when "00001000010010",
                      414 when "00001000010011",
                      413 when "00001000010100",
                      412 when "00001000010101",
                      411 when "00001000010110",
                      411 when "00001000010111",
                      410 when "00001000011000",
                      409 when "00001000011001",
                      408 when "00001000011010",
                      408 when "00001000011011",
                      407 when "00001000011100",
                      406 when "00001000011101",
                      405 when "00001000011110",
                      405 when "00001000011111",
                      404 when "00001000100000",
                      403 when "00001000100001",
                      402 when "00001000100010",
                      402 when "00001000100011",
                      401 when "00001000100100",
                      400 when "00001000100101",
                      400 when "00001000100110",
                      399 when "00001000100111",
                      398 when "00001000101000",
                      397 when "00001000101001",
                      397 when "00001000101010",
                      396 when "00001000101011",
                      395 when "00001000101100",
                      394 when "00001000101101",
                      394 when "00001000101110",
                      393 when "00001000101111",
                      392 when "00001000110000",
                      392 when "00001000110001",
                      391 when "00001000110010",
                      390 when "00001000110011",
                      390 when "00001000110100",
                      389 when "00001000110101",
                      388 when "00001000110110",
                      388 when "00001000110111",
                      387 when "00001000111000",
                      386 when "00001000111001",
                      385 when "00001000111010",
                      385 when "00001000111011",
                      384 when "00001000111100",
                      383 when "00001000111101",
                      383 when "00001000111110",
                      382 when "00001000111111",
                      381 when "00001001000000",
                      381 when "00001001000001",
                      380 when "00001001000010",
                      379 when "00001001000011",
                      379 when "00001001000100",
                      378 when "00001001000101",
                      378 when "00001001000110",
                      377 when "00001001000111",
                      376 when "00001001001000",
                      376 when "00001001001001",
                      375 when "00001001001010",
                      374 when "00001001001011",
                      374 when "00001001001100",
                      373 when "00001001001101",
                      372 when "00001001001110",
                      372 when "00001001001111",
                      371 when "00001001010000",
                      371 when "00001001010001",
                      370 when "00001001010010",
                      369 when "00001001010011",
                      369 when "00001001010100",
                      368 when "00001001010101",
                      367 when "00001001010110",
                      367 when "00001001010111",
                      366 when "00001001011000",
                      366 when "00001001011001",
                      365 when "00001001011010",
                      364 when "00001001011011",
                      364 when "00001001011100",
                      363 when "00001001011101",
                      363 when "00001001011110",
                      362 when "00001001011111",
                      361 when "00001001100000",
                      361 when "00001001100001",
                      360 when "00001001100010",
                      360 when "00001001100011",
                      359 when "00001001100100",
                      358 when "00001001100101",
                      358 when "00001001100110",
                      357 when "00001001100111",
                      357 when "00001001101000",
                      356 when "00001001101001",
                      356 when "00001001101010",
                      355 when "00001001101011",
                      354 when "00001001101100",
                      354 when "00001001101101",
                      353 when "00001001101110",
                      353 when "00001001101111",
                      352 when "00001001110000",
                      352 when "00001001110001",
                      351 when "00001001110010",
                      350 when "00001001110011",
                      350 when "00001001110100",
                      349 when "00001001110101",
                      349 when "00001001110110",
                      348 when "00001001110111",
                      348 when "00001001111000",
                      347 when "00001001111001",
                      347 when "00001001111010",
                      346 when "00001001111011",
                      345 when "00001001111100",
                      345 when "00001001111101",
                      344 when "00001001111110",
                      344 when "00001001111111",
                      343 when "00001010000000",
                      343 when "00001010000001",
                      342 when "00001010000010",
                      342 when "00001010000011",
                      341 when "00001010000100",
                      341 when "00001010000101",
                      340 when "00001010000110",
                      340 when "00001010000111",
                      339 when "00001010001000",
                      339 when "00001010001001",
                      338 when "00001010001010",
                      338 when "00001010001011",
                      337 when "00001010001100",
                      336 when "00001010001101",
                      336 when "00001010001110",
                      335 when "00001010001111",
                      335 when "00001010010000",
                      334 when "00001010010001",
                      334 when "00001010010010",
                      333 when "00001010010011",
                      333 when "00001010010100",
                      332 when "00001010010101",
                      332 when "00001010010110",
                      331 when "00001010010111",
                      331 when "00001010011000",
                      330 when "00001010011001",
                      330 when "00001010011010",
                      329 when "00001010011011",
                      329 when "00001010011100",
                      328 when "00001010011101",
                      328 when "00001010011110",
                      327 when "00001010011111",
                      327 when "00001010100000",
                      326 when "00001010100001",
                      326 when "00001010100010",
                      326 when "00001010100011",
                      325 when "00001010100100",
                      325 when "00001010100101",
                      324 when "00001010100110",
                      324 when "00001010100111",
                      323 when "00001010101000",
                      323 when "00001010101001",
                      322 when "00001010101010",
                      322 when "00001010101011",
                      321 when "00001010101100",
                      321 when "00001010101101",
                      320 when "00001010101110",
                      320 when "00001010101111",
                      319 when "00001010110000",
                      319 when "00001010110001",
                      318 when "00001010110010",
                      318 when "00001010110011",
                      318 when "00001010110100",
                      317 when "00001010110101",
                      317 when "00001010110110",
                      316 when "00001010110111",
                      316 when "00001010111000",
                      315 when "00001010111001",
                      315 when "00001010111010",
                      314 when "00001010111011",
                      314 when "00001010111100",
                      313 when "00001010111101",
                      313 when "00001010111110",
                      313 when "00001010111111",
                      312 when "00001011000000",
                      312 when "00001011000001",
                      311 when "00001011000010",
                      311 when "00001011000011",
                      310 when "00001011000100",
                      310 when "00001011000101",
                      309 when "00001011000110",
                      309 when "00001011000111",
                      309 when "00001011001000",
                      308 when "00001011001001",
                      308 when "00001011001010",
                      307 when "00001011001011",
                      307 when "00001011001100",
                      306 when "00001011001101",
                      306 when "00001011001110",
                      306 when "00001011001111",
                      305 when "00001011010000",
                      305 when "00001011010001",
                      304 when "00001011010010",
                      304 when "00001011010011",
                      303 when "00001011010100",
                      303 when "00001011010101",
                      303 when "00001011010110",
                      302 when "00001011010111",
                      302 when "00001011011000",
                      301 when "00001011011001",
                      301 when "00001011011010",
                      301 when "00001011011011",
                      300 when "00001011011100",
                      300 when "00001011011101",
                      299 when "00001011011110",
                      299 when "00001011011111",
                      299 when "00001011100000",
                      298 when "00001011100001",
                      298 when "00001011100010",
                      297 when "00001011100011",
                      297 when "00001011100100",
                      297 when "00001011100101",
                      296 when "00001011100110",
                      296 when "00001011100111",
                      295 when "00001011101000",
                      295 when "00001011101001",
                      295 when "00001011101010",
                      294 when "00001011101011",
                      294 when "00001011101100",
                      293 when "00001011101101",
                      293 when "00001011101110",
                      293 when "00001011101111",
                      292 when "00001011110000",
                      292 when "00001011110001",
                      291 when "00001011110010",
                      291 when "00001011110011",
                      291 when "00001011110100",
                      290 when "00001011110101",
                      290 when "00001011110110",
                      289 when "00001011110111",
                      289 when "00001011111000",
                      289 when "00001011111001",
                      288 when "00001011111010",
                      288 when "00001011111011",
                      288 when "00001011111100",
                      287 when "00001011111101",
                      287 when "00001011111110",
                      286 when "00001011111111",
                      286 when "00001100000000",
                      286 when "00001100000001",
                      285 when "00001100000010",
                      285 when "00001100000011",
                      285 when "00001100000100",
                      284 when "00001100000101",
                      284 when "00001100000110",
                      284 when "00001100000111",
                      283 when "00001100001000",
                      283 when "00001100001001",
                      282 when "00001100001010",
                      282 when "00001100001011",
                      282 when "00001100001100",
                      281 when "00001100001101",
                      281 when "00001100001110",
                      281 when "00001100001111",
                      280 when "00001100010000",
                      280 when "00001100010001",
                      280 when "00001100010010",
                      279 when "00001100010011",
                      279 when "00001100010100",
                      278 when "00001100010101",
                      278 when "00001100010110",
                      278 when "00001100010111",
                      277 when "00001100011000",
                      277 when "00001100011001",
                      277 when "00001100011010",
                      276 when "00001100011011",
                      276 when "00001100011100",
                      276 when "00001100011101",
                      275 when "00001100011110",
                      275 when "00001100011111",
                      275 when "00001100100000",
                      274 when "00001100100001",
                      274 when "00001100100010",
                      274 when "00001100100011",
                      273 when "00001100100100",
                      273 when "00001100100101",
                      273 when "00001100100110",
                      272 when "00001100100111",
                      272 when "00001100101000",
                      272 when "00001100101001",
                      271 when "00001100101010",
                      271 when "00001100101011",
                      271 when "00001100101100",
                      270 when "00001100101101",
                      270 when "00001100101110",
                      270 when "00001100101111",
                      269 when "00001100110000",
                      269 when "00001100110001",
                      269 when "00001100110010",
                      268 when "00001100110011",
                      268 when "00001100110100",
                      268 when "00001100110101",
                      267 when "00001100110110",
                      267 when "00001100110111",
                      267 when "00001100111000",
                      266 when "00001100111001",
                      266 when "00001100111010",
                      266 when "00001100111011",
                      265 when "00001100111100",
                      265 when "00001100111101",
                      265 when "00001100111110",
                      264 when "00001100111111",
                      264 when "00001101000000",
                      264 when "00001101000001",
                      263 when "00001101000010",
                      263 when "00001101000011",
                      263 when "00001101000100",
                      263 when "00001101000101",
                      262 when "00001101000110",
                      262 when "00001101000111",
                      262 when "00001101001000",
                      261 when "00001101001001",
                      261 when "00001101001010",
                      261 when "00001101001011",
                      260 when "00001101001100",
                      260 when "00001101001101",
                      260 when "00001101001110",
                      259 when "00001101001111",
                      259 when "00001101010000",
                      259 when "00001101010001",
                      259 when "00001101010010",
                      258 when "00001101010011",
                      258 when "00001101010100",
                      258 when "00001101010101",
                      257 when "00001101010110",
                      257 when "00001101010111",
                      257 when "00001101011000",
                      256 when "00001101011001",
                      256 when "00001101011010",
                      256 when "00001101011011",
                      255 when "00001101011100",
                      255 when "00001101011101",
                      255 when "00001101011110",
                      255 when "00001101011111",
                      254 when "00001101100000",
                      254 when "00001101100001",
                      254 when "00001101100010",
                      253 when "00001101100011",
                      253 when "00001101100100",
                      253 when "00001101100101",
                      253 when "00001101100110",
                      252 when "00001101100111",
                      252 when "00001101101000",
                      252 when "00001101101001",
                      251 when "00001101101010",
                      251 when "00001101101011",
                      251 when "00001101101100",
                      251 when "00001101101101",
                      250 when "00001101101110",
                      250 when "00001101101111",
                      250 when "00001101110000",
                      249 when "00001101110001",
                      249 when "00001101110010",
                      249 when "00001101110011",
                      249 when "00001101110100",
                      248 when "00001101110101",
                      248 when "00001101110110",
                      248 when "00001101110111",
                      247 when "00001101111000",
                      247 when "00001101111001",
                      247 when "00001101111010",
                      247 when "00001101111011",
                      246 when "00001101111100",
                      246 when "00001101111101",
                      246 when "00001101111110",
                      246 when "00001101111111",
                      245 when "00001110000000",
                      245 when "00001110000001",
                      245 when "00001110000010",
                      244 when "00001110000011",
                      244 when "00001110000100",
                      244 when "00001110000101",
                      244 when "00001110000110",
                      243 when "00001110000111",
                      243 when "00001110001000",
                      243 when "00001110001001",
                      243 when "00001110001010",
                      242 when "00001110001011",
                      242 when "00001110001100",
                      242 when "00001110001101",
                      241 when "00001110001110",
                      241 when "00001110001111",
                      241 when "00001110010000",
                      241 when "00001110010001",
                      240 when "00001110010010",
                      240 when "00001110010011",
                      240 when "00001110010100",
                      240 when "00001110010101",
                      239 when "00001110010110",
                      239 when "00001110010111",
                      239 when "00001110011000",
                      239 when "00001110011001",
                      238 when "00001110011010",
                      238 when "00001110011011",
                      238 when "00001110011100",
                      238 when "00001110011101",
                      237 when "00001110011110",
                      237 when "00001110011111",
                      237 when "00001110100000",
                      237 when "00001110100001",
                      236 when "00001110100010",
                      236 when "00001110100011",
                      236 when "00001110100100",
                      236 when "00001110100101",
                      235 when "00001110100110",
                      235 when "00001110100111",
                      235 when "00001110101000",
                      235 when "00001110101001",
                      234 when "00001110101010",
                      234 when "00001110101011",
                      234 when "00001110101100",
                      234 when "00001110101101",
                      233 when "00001110101110",
                      233 when "00001110101111",
                      233 when "00001110110000",
                      233 when "00001110110001",
                      232 when "00001110110010",
                      232 when "00001110110011",
                      232 when "00001110110100",
                      232 when "00001110110101",
                      231 when "00001110110110",
                      231 when "00001110110111",
                      231 when "00001110111000",
                      231 when "00001110111001",
                      230 when "00001110111010",
                      230 when "00001110111011",
                      230 when "00001110111100",
                      230 when "00001110111101",
                      229 when "00001110111110",
                      229 when "00001110111111",
                      229 when "00001111000000",
                      229 when "00001111000001",
                      228 when "00001111000010",
                      228 when "00001111000011",
                      228 when "00001111000100",
                      228 when "00001111000101",
                      227 when "00001111000110",
                      227 when "00001111000111",
                      227 when "00001111001000",
                      227 when "00001111001001",
                      227 when "00001111001010",
                      226 when "00001111001011",
                      226 when "00001111001100",
                      226 when "00001111001101",
                      226 when "00001111001110",
                      225 when "00001111001111",
                      225 when "00001111010000",
                      225 when "00001111010001",
                      225 when "00001111010010",
                      224 when "00001111010011",
                      224 when "00001111010100",
                      224 when "00001111010101",
                      224 when "00001111010110",
                      224 when "00001111010111",
                      223 when "00001111011000",
                      223 when "00001111011001",
                      223 when "00001111011010",
                      223 when "00001111011011",
                      222 when "00001111011100",
                      222 when "00001111011101",
                      222 when "00001111011110",
                      222 when "00001111011111",
                      221 when "00001111100000",
                      221 when "00001111100001",
                      221 when "00001111100010",
                      221 when "00001111100011",
                      221 when "00001111100100",
                      220 when "00001111100101",
                      220 when "00001111100110",
                      220 when "00001111100111",
                      220 when "00001111101000",
                      220 when "00001111101001",
                      219 when "00001111101010",
                      219 when "00001111101011",
                      219 when "00001111101100",
                      219 when "00001111101101",
                      218 when "00001111101110",
                      218 when "00001111101111",
                      218 when "00001111110000",
                      218 when "00001111110001",
                      218 when "00001111110010",
                      217 when "00001111110011",
                      217 when "00001111110100",
                      217 when "00001111110101",
                      217 when "00001111110110",
                      216 when "00001111110111",
                      216 when "00001111111000",
                      216 when "00001111111001",
                      216 when "00001111111010",
                      216 when "00001111111011",
                      215 when "00001111111100",
                      215 when "00001111111101",
                      215 when "00001111111110",
                      215 when "00001111111111",
                      215 when "00010000000000",
                      214 when "00010000000001",
                      214 when "00010000000010",
                      214 when "00010000000011",
                      214 when "00010000000100",
                      214 when "00010000000101",
                      213 when "00010000000110",
                      213 when "00010000000111",
                      213 when "00010000001000",
                      213 when "00010000001001",
                      213 when "00010000001010",
                      212 when "00010000001011",
                      212 when "00010000001100",
                      212 when "00010000001101",
                      212 when "00010000001110",
                      211 when "00010000001111",
                      211 when "00010000010000",
                      211 when "00010000010001",
                      211 when "00010000010010",
                      211 when "00010000010011",
                      210 when "00010000010100",
                      210 when "00010000010101",
                      210 when "00010000010110",
                      210 when "00010000010111",
                      210 when "00010000011000",
                      209 when "00010000011001",
                      209 when "00010000011010",
                      209 when "00010000011011",
                      209 when "00010000011100",
                      209 when "00010000011101",
                      208 when "00010000011110",
                      208 when "00010000011111",
                      208 when "00010000100000",
                      208 when "00010000100001",
                      208 when "00010000100010",
                      207 when "00010000100011",
                      207 when "00010000100100",
                      207 when "00010000100101",
                      207 when "00010000100110",
                      207 when "00010000100111",
                      207 when "00010000101000",
                      206 when "00010000101001",
                      206 when "00010000101010",
                      206 when "00010000101011",
                      206 when "00010000101100",
                      206 when "00010000101101",
                      205 when "00010000101110",
                      205 when "00010000101111",
                      205 when "00010000110000",
                      205 when "00010000110001",
                      205 when "00010000110010",
                      204 when "00010000110011",
                      204 when "00010000110100",
                      204 when "00010000110101",
                      204 when "00010000110110",
                      204 when "00010000110111",
                      203 when "00010000111000",
                      203 when "00010000111001",
                      203 when "00010000111010",
                      203 when "00010000111011",
                      203 when "00010000111100",
                      203 when "00010000111101",
                      202 when "00010000111110",
                      202 when "00010000111111",
                      202 when "00010001000000",
                      202 when "00010001000001",
                      202 when "00010001000010",
                      201 when "00010001000011",
                      201 when "00010001000100",
                      201 when "00010001000101",
                      201 when "00010001000110",
                      201 when "00010001000111",
                      200 when "00010001001000",
                      200 when "00010001001001",
                      200 when "00010001001010",
                      200 when "00010001001011",
                      200 when "00010001001100",
                      200 when "00010001001101",
                      199 when "00010001001110",
                      199 when "00010001001111",
                      199 when "00010001010000",
                      199 when "00010001010001",
                      199 when "00010001010010",
                      198 when "00010001010011",
                      198 when "00010001010100",
                      198 when "00010001010101",
                      198 when "00010001010110",
                      198 when "00010001010111",
                      198 when "00010001011000",
                      197 when "00010001011001",
                      197 when "00010001011010",
                      197 when "00010001011011",
                      197 when "00010001011100",
                      197 when "00010001011101",
                      197 when "00010001011110",
                      196 when "00010001011111",
                      196 when "00010001100000",
                      196 when "00010001100001",
                      196 when "00010001100010",
                      196 when "00010001100011",
                      195 when "00010001100100",
                      195 when "00010001100101",
                      195 when "00010001100110",
                      195 when "00010001100111",
                      195 when "00010001101000",
                      195 when "00010001101001",
                      194 when "00010001101010",
                      194 when "00010001101011",
                      194 when "00010001101100",
                      194 when "00010001101101",
                      194 when "00010001101110",
                      194 when "00010001101111",
                      193 when "00010001110000",
                      193 when "00010001110001",
                      193 when "00010001110010",
                      193 when "00010001110011",
                      193 when "00010001110100",
                      193 when "00010001110101",
                      192 when "00010001110110",
                      192 when "00010001110111",
                      192 when "00010001111000",
                      192 when "00010001111001",
                      192 when "00010001111010",
                      192 when "00010001111011",
                      191 when "00010001111100",
                      191 when "00010001111101",
                      191 when "00010001111110",
                      191 when "00010001111111",
                      191 when "00010010000000",
                      191 when "00010010000001",
                      190 when "00010010000010",
                      190 when "00010010000011",
                      190 when "00010010000100",
                      190 when "00010010000101",
                      190 when "00010010000110",
                      190 when "00010010000111",
                      189 when "00010010001000",
                      189 when "00010010001001",
                      189 when "00010010001010",
                      189 when "00010010001011",
                      189 when "00010010001100",
                      189 when "00010010001101",
                      188 when "00010010001110",
                      188 when "00010010001111",
                      188 when "00010010010000",
                      188 when "00010010010001",
                      188 when "00010010010010",
                      188 when "00010010010011",
                      187 when "00010010010100",
                      187 when "00010010010101",
                      187 when "00010010010110",
                      187 when "00010010010111",
                      187 when "00010010011000",
                      187 when "00010010011001",
                      187 when "00010010011010",
                      186 when "00010010011011",
                      186 when "00010010011100",
                      186 when "00010010011101",
                      186 when "00010010011110",
                      186 when "00010010011111",
                      186 when "00010010100000",
                      185 when "00010010100001",
                      185 when "00010010100010",
                      185 when "00010010100011",
                      185 when "00010010100100",
                      185 when "00010010100101",
                      185 when "00010010100110",
                      184 when "00010010100111",
                      184 when "00010010101000",
                      184 when "00010010101001",
                      184 when "00010010101010",
                      184 when "00010010101011",
                      184 when "00010010101100",
                      184 when "00010010101101",
                      183 when "00010010101110",
                      183 when "00010010101111",
                      183 when "00010010110000",
                      183 when "00010010110001",
                      183 when "00010010110010",
                      183 when "00010010110011",
                      182 when "00010010110100",
                      182 when "00010010110101",
                      182 when "00010010110110",
                      182 when "00010010110111",
                      182 when "00010010111000",
                      182 when "00010010111001",
                      182 when "00010010111010",
                      181 when "00010010111011",
                      181 when "00010010111100",
                      181 when "00010010111101",
                      181 when "00010010111110",
                      181 when "00010010111111",
                      181 when "00010011000000",
                      181 when "00010011000001",
                      180 when "00010011000010",
                      180 when "00010011000011",
                      180 when "00010011000100",
                      180 when "00010011000101",
                      180 when "00010011000110",
                      180 when "00010011000111",
                      180 when "00010011001000",
                      179 when "00010011001001",
                      179 when "00010011001010",
                      179 when "00010011001011",
                      179 when "00010011001100",
                      179 when "00010011001101",
                      179 when "00010011001110",
                      178 when "00010011001111",
                      178 when "00010011010000",
                      178 when "00010011010001",
                      178 when "00010011010010",
                      178 when "00010011010011",
                      178 when "00010011010100",
                      178 when "00010011010101",
                      177 when "00010011010110",
                      177 when "00010011010111",
                      177 when "00010011011000",
                      177 when "00010011011001",
                      177 when "00010011011010",
                      177 when "00010011011011",
                      177 when "00010011011100",
                      176 when "00010011011101",
                      176 when "00010011011110",
                      176 when "00010011011111",
                      176 when "00010011100000",
                      176 when "00010011100001",
                      176 when "00010011100010",
                      176 when "00010011100011",
                      176 when "00010011100100",
                      175 when "00010011100101",
                      175 when "00010011100110",
                      175 when "00010011100111",
                      175 when "00010011101000",
                      175 when "00010011101001",
                      175 when "00010011101010",
                      175 when "00010011101011",
                      174 when "00010011101100",
                      174 when "00010011101101",
                      174 when "00010011101110",
                      174 when "00010011101111",
                      174 when "00010011110000",
                      174 when "00010011110001",
                      174 when "00010011110010",
                      173 when "00010011110011",
                      173 when "00010011110100",
                      173 when "00010011110101",
                      173 when "00010011110110",
                      173 when "00010011110111",
                      173 when "00010011111000",
                      173 when "00010011111001",
                      172 when "00010011111010",
                      172 when "00010011111011",
                      172 when "00010011111100",
                      172 when "00010011111101",
                      172 when "00010011111110",
                      172 when "00010011111111",
                      172 when "00010100000000",
                      172 when "00010100000001",
                      171 when "00010100000010",
                      171 when "00010100000011",
                      171 when "00010100000100",
                      171 when "00010100000101",
                      171 when "00010100000110",
                      171 when "00010100000111",
                      171 when "00010100001000",
                      170 when "00010100001001",
                      170 when "00010100001010",
                      170 when "00010100001011",
                      170 when "00010100001100",
                      170 when "00010100001101",
                      170 when "00010100001110",
                      170 when "00010100001111",
                      170 when "00010100010000",
                      169 when "00010100010001",
                      169 when "00010100010010",
                      169 when "00010100010011",
                      169 when "00010100010100",
                      169 when "00010100010101",
                      169 when "00010100010110",
                      169 when "00010100010111",
                      169 when "00010100011000",
                      168 when "00010100011001",
                      168 when "00010100011010",
                      168 when "00010100011011",
                      168 when "00010100011100",
                      168 when "00010100011101",
                      168 when "00010100011110",
                      168 when "00010100011111",
                      167 when "00010100100000",
                      167 when "00010100100001",
                      167 when "00010100100010",
                      167 when "00010100100011",
                      167 when "00010100100100",
                      167 when "00010100100101",
                      167 when "00010100100110",
                      167 when "00010100100111",
                      166 when "00010100101000",
                      166 when "00010100101001",
                      166 when "00010100101010",
                      166 when "00010100101011",
                      166 when "00010100101100",
                      166 when "00010100101101",
                      166 when "00010100101110",
                      166 when "00010100101111",
                      165 when "00010100110000",
                      165 when "00010100110001",
                      165 when "00010100110010",
                      165 when "00010100110011",
                      165 when "00010100110100",
                      165 when "00010100110101",
                      165 when "00010100110110",
                      165 when "00010100110111",
                      164 when "00010100111000",
                      164 when "00010100111001",
                      164 when "00010100111010",
                      164 when "00010100111011",
                      164 when "00010100111100",
                      164 when "00010100111101",
                      164 when "00010100111110",
                      164 when "00010100111111",
                      163 when "00010101000000",
                      163 when "00010101000001",
                      163 when "00010101000010",
                      163 when "00010101000011",
                      163 when "00010101000100",
                      163 when "00010101000101",
                      163 when "00010101000110",
                      163 when "00010101000111",
                      163 when "00010101001000",
                      162 when "00010101001001",
                      162 when "00010101001010",
                      162 when "00010101001011",
                      162 when "00010101001100",
                      162 when "00010101001101",
                      162 when "00010101001110",
                      162 when "00010101001111",
                      162 when "00010101010000",
                      161 when "00010101010001",
                      161 when "00010101010010",
                      161 when "00010101010011",
                      161 when "00010101010100",
                      161 when "00010101010101",
                      161 when "00010101010110",
                      161 when "00010101010111",
                      161 when "00010101011000",
                      161 when "00010101011001",
                      160 when "00010101011010",
                      160 when "00010101011011",
                      160 when "00010101011100",
                      160 when "00010101011101",
                      160 when "00010101011110",
                      160 when "00010101011111",
                      160 when "00010101100000",
                      160 when "00010101100001",
                      159 when "00010101100010",
                      159 when "00010101100011",
                      159 when "00010101100100",
                      159 when "00010101100101",
                      159 when "00010101100110",
                      159 when "00010101100111",
                      159 when "00010101101000",
                      159 when "00010101101001",
                      159 when "00010101101010",
                      158 when "00010101101011",
                      158 when "00010101101100",
                      158 when "00010101101101",
                      158 when "00010101101110",
                      158 when "00010101101111",
                      158 when "00010101110000",
                      158 when "00010101110001",
                      158 when "00010101110010",
                      158 when "00010101110011",
                      157 when "00010101110100",
                      157 when "00010101110101",
                      157 when "00010101110110",
                      157 when "00010101110111",
                      157 when "00010101111000",
                      157 when "00010101111001",
                      157 when "00010101111010",
                      157 when "00010101111011",
                      157 when "00010101111100",
                      156 when "00010101111101",
                      156 when "00010101111110",
                      156 when "00010101111111",
                      156 when "00010110000000",
                      156 when "00010110000001",
                      156 when "00010110000010",
                      156 when "00010110000011",
                      156 when "00010110000100",
                      156 when "00010110000101",
                      155 when "00010110000110",
                      155 when "00010110000111",
                      155 when "00010110001000",
                      155 when "00010110001001",
                      155 when "00010110001010",
                      155 when "00010110001011",
                      155 when "00010110001100",
                      155 when "00010110001101",
                      155 when "00010110001110",
                      154 when "00010110001111",
                      154 when "00010110010000",
                      154 when "00010110010001",
                      154 when "00010110010010",
                      154 when "00010110010011",
                      154 when "00010110010100",
                      154 when "00010110010101",
                      154 when "00010110010110",
                      154 when "00010110010111",
                      153 when "00010110011000",
                      153 when "00010110011001",
                      153 when "00010110011010",
                      153 when "00010110011011",
                      153 when "00010110011100",
                      153 when "00010110011101",
                      153 when "00010110011110",
                      153 when "00010110011111",
                      153 when "00010110100000",
                      152 when "00010110100001",
                      152 when "00010110100010",
                      152 when "00010110100011",
                      152 when "00010110100100",
                      152 when "00010110100101",
                      152 when "00010110100110",
                      152 when "00010110100111",
                      152 when "00010110101000",
                      152 when "00010110101001",
                      152 when "00010110101010",
                      151 when "00010110101011",
                      151 when "00010110101100",
                      151 when "00010110101101",
                      151 when "00010110101110",
                      151 when "00010110101111",
                      151 when "00010110110000",
                      151 when "00010110110001",
                      151 when "00010110110010",
                      151 when "00010110110011",
                      150 when "00010110110100",
                      150 when "00010110110101",
                      150 when "00010110110110",
                      150 when "00010110110111",
                      150 when "00010110111000",
                      150 when "00010110111001",
                      150 when "00010110111010",
                      150 when "00010110111011",
                      150 when "00010110111100",
                      150 when "00010110111101",
                      149 when "00010110111110",
                      149 when "00010110111111",
                      149 when "00010111000000",
                      149 when "00010111000001",
                      149 when "00010111000010",
                      149 when "00010111000011",
                      149 when "00010111000100",
                      149 when "00010111000101",
                      149 when "00010111000110",
                      149 when "00010111000111",
                      148 when "00010111001000",
                      148 when "00010111001001",
                      148 when "00010111001010",
                      148 when "00010111001011",
                      148 when "00010111001100",
                      148 when "00010111001101",
                      148 when "00010111001110",
                      148 when "00010111001111",
                      148 when "00010111010000",
                      148 when "00010111010001",
                      147 when "00010111010010",
                      147 when "00010111010011",
                      147 when "00010111010100",
                      147 when "00010111010101",
                      147 when "00010111010110",
                      147 when "00010111010111",
                      147 when "00010111011000",
                      147 when "00010111011001",
                      147 when "00010111011010",
                      147 when "00010111011011",
                      146 when "00010111011100",
                      146 when "00010111011101",
                      146 when "00010111011110",
                      146 when "00010111011111",
                      146 when "00010111100000",
                      146 when "00010111100001",
                      146 when "00010111100010",
                      146 when "00010111100011",
                      146 when "00010111100100",
                      146 when "00010111100101",
                      146 when "00010111100110",
                      145 when "00010111100111",
                      145 when "00010111101000",
                      145 when "00010111101001",
                      145 when "00010111101010",
                      145 when "00010111101011",
                      145 when "00010111101100",
                      145 when "00010111101101",
                      145 when "00010111101110",
                      145 when "00010111101111",
                      145 when "00010111110000",
                      144 when "00010111110001",
                      144 when "00010111110010",
                      144 when "00010111110011",
                      144 when "00010111110100",
                      144 when "00010111110101",
                      144 when "00010111110110",
                      144 when "00010111110111",
                      144 when "00010111111000",
                      144 when "00010111111001",
                      144 when "00010111111010",
                      144 when "00010111111011",
                      143 when "00010111111100",
                      143 when "00010111111101",
                      143 when "00010111111110",
                      143 when "00010111111111",
                      143 when "00011000000000",
                      143 when "00011000000001",
                      143 when "00011000000010",
                      143 when "00011000000011",
                      143 when "00011000000100",
                      143 when "00011000000101",
                      142 when "00011000000110",
                      142 when "00011000000111",
                      142 when "00011000001000",
                      142 when "00011000001001",
                      142 when "00011000001010",
                      142 when "00011000001011",
                      142 when "00011000001100",
                      142 when "00011000001101",
                      142 when "00011000001110",
                      142 when "00011000001111",
                      142 when "00011000010000",
                      141 when "00011000010001",
                      141 when "00011000010010",
                      141 when "00011000010011",
                      141 when "00011000010100",
                      141 when "00011000010101",
                      141 when "00011000010110",
                      141 when "00011000010111",
                      141 when "00011000011000",
                      141 when "00011000011001",
                      141 when "00011000011010",
                      141 when "00011000011011",
                      140 when "00011000011100",
                      140 when "00011000011101",
                      140 when "00011000011110",
                      140 when "00011000011111",
                      140 when "00011000100000",
                      140 when "00011000100001",
                      140 when "00011000100010",
                      140 when "00011000100011",
                      140 when "00011000100100",
                      140 when "00011000100101",
                      140 when "00011000100110",
                      140 when "00011000100111",
                      139 when "00011000101000",
                      139 when "00011000101001",
                      139 when "00011000101010",
                      139 when "00011000101011",
                      139 when "00011000101100",
                      139 when "00011000101101",
                      139 when "00011000101110",
                      139 when "00011000101111",
                      139 when "00011000110000",
                      139 when "00011000110001",
                      139 when "00011000110010",
                      138 when "00011000110011",
                      138 when "00011000110100",
                      138 when "00011000110101",
                      138 when "00011000110110",
                      138 when "00011000110111",
                      138 when "00011000111000",
                      138 when "00011000111001",
                      138 when "00011000111010",
                      138 when "00011000111011",
                      138 when "00011000111100",
                      138 when "00011000111101",
                      138 when "00011000111110",
                      137 when "00011000111111",
                      137 when "00011001000000",
                      137 when "00011001000001",
                      137 when "00011001000010",
                      137 when "00011001000011",
                      137 when "00011001000100",
                      137 when "00011001000101",
                      137 when "00011001000110",
                      137 when "00011001000111",
                      137 when "00011001001000",
                      137 when "00011001001001",
                      136 when "00011001001010",
                      136 when "00011001001011",
                      136 when "00011001001100",
                      136 when "00011001001101",
                      136 when "00011001001110",
                      136 when "00011001001111",
                      136 when "00011001010000",
                      136 when "00011001010001",
                      136 when "00011001010010",
                      136 when "00011001010011",
                      136 when "00011001010100",
                      136 when "00011001010101",
                      135 when "00011001010110",
                      135 when "00011001010111",
                      135 when "00011001011000",
                      135 when "00011001011001",
                      135 when "00011001011010",
                      135 when "00011001011011",
                      135 when "00011001011100",
                      135 when "00011001011101",
                      135 when "00011001011110",
                      135 when "00011001011111",
                      135 when "00011001100000",
                      135 when "00011001100001",
                      134 when "00011001100010",
                      134 when "00011001100011",
                      134 when "00011001100100",
                      134 when "00011001100101",
                      134 when "00011001100110",
                      134 when "00011001100111",
                      134 when "00011001101000",
                      134 when "00011001101001",
                      134 when "00011001101010",
                      134 when "00011001101011",
                      134 when "00011001101100",
                      134 when "00011001101101",
                      133 when "00011001101110",
                      133 when "00011001101111",
                      133 when "00011001110000",
                      133 when "00011001110001",
                      133 when "00011001110010",
                      133 when "00011001110011",
                      133 when "00011001110100",
                      133 when "00011001110101",
                      133 when "00011001110110",
                      133 when "00011001110111",
                      133 when "00011001111000",
                      133 when "00011001111001",
                      133 when "00011001111010",
                      132 when "00011001111011",
                      132 when "00011001111100",
                      132 when "00011001111101",
                      132 when "00011001111110",
                      132 when "00011001111111",
                      132 when "00011010000000",
                      132 when "00011010000001",
                      132 when "00011010000010",
                      132 when "00011010000011",
                      132 when "00011010000100",
                      132 when "00011010000101",
                      132 when "00011010000110",
                      131 when "00011010000111",
                      131 when "00011010001000",
                      131 when "00011010001001",
                      131 when "00011010001010",
                      131 when "00011010001011",
                      131 when "00011010001100",
                      131 when "00011010001101",
                      131 when "00011010001110",
                      131 when "00011010001111",
                      131 when "00011010010000",
                      131 when "00011010010001",
                      131 when "00011010010010",
                      131 when "00011010010011",
                      130 when "00011010010100",
                      130 when "00011010010101",
                      130 when "00011010010110",
                      130 when "00011010010111",
                      130 when "00011010011000",
                      130 when "00011010011001",
                      130 when "00011010011010",
                      130 when "00011010011011",
                      130 when "00011010011100",
                      130 when "00011010011101",
                      130 when "00011010011110",
                      130 when "00011010011111",
                      130 when "00011010100000",
                      129 when "00011010100001",
                      129 when "00011010100010",
                      129 when "00011010100011",
                      129 when "00011010100100",
                      129 when "00011010100101",
                      129 when "00011010100110",
                      129 when "00011010100111",
                      129 when "00011010101000",
                      129 when "00011010101001",
                      129 when "00011010101010",
                      129 when "00011010101011",
                      129 when "00011010101100",
                      129 when "00011010101101",
                      128 when "00011010101110",
                      128 when "00011010101111",
                      128 when "00011010110000",
                      128 when "00011010110001",
                      128 when "00011010110010",
                      128 when "00011010110011",
                      128 when "00011010110100",
                      128 when "00011010110101",
                      128 when "00011010110110",
                      128 when "00011010110111",
                      128 when "00011010111000",
                      128 when "00011010111001",
                      128 when "00011010111010",
                      128 when "00011010111011",
                      127 when "00011010111100",
                      127 when "00011010111101",
                      127 when "00011010111110",
                      127 when "00011010111111",
                      127 when "00011011000000",
                      127 when "00011011000001",
                      127 when "00011011000010",
                      127 when "00011011000011",
                      127 when "00011011000100",
                      127 when "00011011000101",
                      127 when "00011011000110",
                      127 when "00011011000111",
                      127 when "00011011001000",
                      126 when "00011011001001",
                      126 when "00011011001010",
                      126 when "00011011001011",
                      126 when "00011011001100",
                      126 when "00011011001101",
                      126 when "00011011001110",
                      126 when "00011011001111",
                      126 when "00011011010000",
                      126 when "00011011010001",
                      126 when "00011011010010",
                      126 when "00011011010011",
                      126 when "00011011010100",
                      126 when "00011011010101",
                      126 when "00011011010110",
                      125 when "00011011010111",
                      125 when "00011011011000",
                      125 when "00011011011001",
                      125 when "00011011011010",
                      125 when "00011011011011",
                      125 when "00011011011100",
                      125 when "00011011011101",
                      125 when "00011011011110",
                      125 when "00011011011111",
                      125 when "00011011100000",
                      125 when "00011011100001",
                      125 when "00011011100010",
                      125 when "00011011100011",
                      125 when "00011011100100",
                      124 when "00011011100101",
                      124 when "00011011100110",
                      124 when "00011011100111",
                      124 when "00011011101000",
                      124 when "00011011101001",
                      124 when "00011011101010",
                      124 when "00011011101011",
                      124 when "00011011101100",
                      124 when "00011011101101",
                      124 when "00011011101110",
                      124 when "00011011101111",
                      124 when "00011011110000",
                      124 when "00011011110001",
                      124 when "00011011110010",
                      124 when "00011011110011",
                      123 when "00011011110100",
                      123 when "00011011110101",
                      123 when "00011011110110",
                      123 when "00011011110111",
                      123 when "00011011111000",
                      123 when "00011011111001",
                      123 when "00011011111010",
                      123 when "00011011111011",
                      123 when "00011011111100",
                      123 when "00011011111101",
                      123 when "00011011111110",
                      123 when "00011011111111",
                      123 when "00011100000000",
                      123 when "00011100000001",
                      122 when "00011100000010",
                      122 when "00011100000011",
                      122 when "00011100000100",
                      122 when "00011100000101",
                      122 when "00011100000110",
                      122 when "00011100000111",
                      122 when "00011100001000",
                      122 when "00011100001001",
                      122 when "00011100001010",
                      122 when "00011100001011",
                      122 when "00011100001100",
                      122 when "00011100001101",
                      122 when "00011100001110",
                      122 when "00011100001111",
                      122 when "00011100010000",
                      121 when "00011100010001",
                      121 when "00011100010010",
                      121 when "00011100010011",
                      121 when "00011100010100",
                      121 when "00011100010101",
                      121 when "00011100010110",
                      121 when "00011100010111",
                      121 when "00011100011000",
                      121 when "00011100011001",
                      121 when "00011100011010",
                      121 when "00011100011011",
                      121 when "00011100011100",
                      121 when "00011100011101",
                      121 when "00011100011110",
                      121 when "00011100011111",
                      120 when "00011100100000",
                      120 when "00011100100001",
                      120 when "00011100100010",
                      120 when "00011100100011",
                      120 when "00011100100100",
                      120 when "00011100100101",
                      120 when "00011100100110",
                      120 when "00011100100111",
                      120 when "00011100101000",
                      120 when "00011100101001",
                      120 when "00011100101010",
                      120 when "00011100101011",
                      120 when "00011100101100",
                      120 when "00011100101101",
                      120 when "00011100101110",
                      119 when "00011100101111",
                      119 when "00011100110000",
                      119 when "00011100110001",
                      119 when "00011100110010",
                      119 when "00011100110011",
                      119 when "00011100110100",
                      119 when "00011100110101",
                      119 when "00011100110110",
                      119 when "00011100110111",
                      119 when "00011100111000",
                      119 when "00011100111001",
                      119 when "00011100111010",
                      119 when "00011100111011",
                      119 when "00011100111100",
                      119 when "00011100111101",
                      119 when "00011100111110",
                      118 when "00011100111111",
                      118 when "00011101000000",
                      118 when "00011101000001",
                      118 when "00011101000010",
                      118 when "00011101000011",
                      118 when "00011101000100",
                      118 when "00011101000101",
                      118 when "00011101000110",
                      118 when "00011101000111",
                      118 when "00011101001000",
                      118 when "00011101001001",
                      118 when "00011101001010",
                      118 when "00011101001011",
                      118 when "00011101001100",
                      118 when "00011101001101",
                      118 when "00011101001110",
                      117 when "00011101001111",
                      117 when "00011101010000",
                      117 when "00011101010001",
                      117 when "00011101010010",
                      117 when "00011101010011",
                      117 when "00011101010100",
                      117 when "00011101010101",
                      117 when "00011101010110",
                      117 when "00011101010111",
                      117 when "00011101011000",
                      117 when "00011101011001",
                      117 when "00011101011010",
                      117 when "00011101011011",
                      117 when "00011101011100",
                      117 when "00011101011101",
                      117 when "00011101011110",
                      116 when "00011101011111",
                      116 when "00011101100000",
                      116 when "00011101100001",
                      116 when "00011101100010",
                      116 when "00011101100011",
                      116 when "00011101100100",
                      116 when "00011101100101",
                      116 when "00011101100110",
                      116 when "00011101100111",
                      116 when "00011101101000",
                      116 when "00011101101001",
                      116 when "00011101101010",
                      116 when "00011101101011",
                      116 when "00011101101100",
                      116 when "00011101101101",
                      116 when "00011101101110",
                      115 when "00011101101111",
                      115 when "00011101110000",
                      115 when "00011101110001",
                      115 when "00011101110010",
                      115 when "00011101110011",
                      115 when "00011101110100",
                      115 when "00011101110101",
                      115 when "00011101110110",
                      115 when "00011101110111",
                      115 when "00011101111000",
                      115 when "00011101111001",
                      115 when "00011101111010",
                      115 when "00011101111011",
                      115 when "00011101111100",
                      115 when "00011101111101",
                      115 when "00011101111110",
                      115 when "00011101111111",
                      114 when "00011110000000",
                      114 when "00011110000001",
                      114 when "00011110000010",
                      114 when "00011110000011",
                      114 when "00011110000100",
                      114 when "00011110000101",
                      114 when "00011110000110",
                      114 when "00011110000111",
                      114 when "00011110001000",
                      114 when "00011110001001",
                      114 when "00011110001010",
                      114 when "00011110001011",
                      114 when "00011110001100",
                      114 when "00011110001101",
                      114 when "00011110001110",
                      114 when "00011110001111",
                      113 when "00011110010000",
                      113 when "00011110010001",
                      113 when "00011110010010",
                      113 when "00011110010011",
                      113 when "00011110010100",
                      113 when "00011110010101",
                      113 when "00011110010110",
                      113 when "00011110010111",
                      113 when "00011110011000",
                      113 when "00011110011001",
                      113 when "00011110011010",
                      113 when "00011110011011",
                      113 when "00011110011100",
                      113 when "00011110011101",
                      113 when "00011110011110",
                      113 when "00011110011111",
                      113 when "00011110100000",
                      113 when "00011110100001",
                      112 when "00011110100010",
                      112 when "00011110100011",
                      112 when "00011110100100",
                      112 when "00011110100101",
                      112 when "00011110100110",
                      112 when "00011110100111",
                      112 when "00011110101000",
                      112 when "00011110101001",
                      112 when "00011110101010",
                      112 when "00011110101011",
                      112 when "00011110101100",
                      112 when "00011110101101",
                      112 when "00011110101110",
                      112 when "00011110101111",
                      112 when "00011110110000",
                      112 when "00011110110001",
                      112 when "00011110110010",
                      111 when "00011110110011",
                      111 when "00011110110100",
                      111 when "00011110110101",
                      111 when "00011110110110",
                      111 when "00011110110111",
                      111 when "00011110111000",
                      111 when "00011110111001",
                      111 when "00011110111010",
                      111 when "00011110111011",
                      111 when "00011110111100",
                      111 when "00011110111101",
                      111 when "00011110111110",
                      111 when "00011110111111",
                      111 when "00011111000000",
                      111 when "00011111000001",
                      111 when "00011111000010",
                      111 when "00011111000011",
                      111 when "00011111000100",
                      110 when "00011111000101",
                      110 when "00011111000110",
                      110 when "00011111000111",
                      110 when "00011111001000",
                      110 when "00011111001001",
                      110 when "00011111001010",
                      110 when "00011111001011",
                      110 when "00011111001100",
                      110 when "00011111001101",
                      110 when "00011111001110",
                      110 when "00011111001111",
                      110 when "00011111010000",
                      110 when "00011111010001",
                      110 when "00011111010010",
                      110 when "00011111010011",
                      110 when "00011111010100",
                      110 when "00011111010101",
                      110 when "00011111010110",
                      109 when "00011111010111",
                      109 when "00011111011000",
                      109 when "00011111011001",
                      109 when "00011111011010",
                      109 when "00011111011011",
                      109 when "00011111011100",
                      109 when "00011111011101",
                      109 when "00011111011110",
                      109 when "00011111011111",
                      109 when "00011111100000",
                      109 when "00011111100001",
                      109 when "00011111100010",
                      109 when "00011111100011",
                      109 when "00011111100100",
                      109 when "00011111100101",
                      109 when "00011111100110",
                      109 when "00011111100111",
                      109 when "00011111101000",
                      109 when "00011111101001",
                      108 when "00011111101010",
                      108 when "00011111101011",
                      108 when "00011111101100",
                      108 when "00011111101101",
                      108 when "00011111101110",
                      108 when "00011111101111",
                      108 when "00011111110000",
                      108 when "00011111110001",
                      108 when "00011111110010",
                      108 when "00011111110011",
                      108 when "00011111110100",
                      108 when "00011111110101",
                      108 when "00011111110110",
                      108 when "00011111110111",
                      108 when "00011111111000",
                      108 when "00011111111001",
                      108 when "00011111111010",
                      108 when "00011111111011",
                      107 when "00011111111100",
                      107 when "00011111111101",
                      107 when "00011111111110",
                      107 when "00011111111111",
                      107 when "00100000000000",
                      107 when "00100000000001",
                      107 when "00100000000010",
                      107 when "00100000000011",
                      107 when "00100000000100",
                      107 when "00100000000101",
                      107 when "00100000000110",
                      107 when "00100000000111",
                      107 when "00100000001000",
                      107 when "00100000001001",
                      107 when "00100000001010",
                      107 when "00100000001011",
                      107 when "00100000001100",
                      107 when "00100000001101",
                      107 when "00100000001110",
                      107 when "00100000001111",
                      106 when "00100000010000",
                      106 when "00100000010001",
                      106 when "00100000010010",
                      106 when "00100000010011",
                      106 when "00100000010100",
                      106 when "00100000010101",
                      106 when "00100000010110",
                      106 when "00100000010111",
                      106 when "00100000011000",
                      106 when "00100000011001",
                      106 when "00100000011010",
                      106 when "00100000011011",
                      106 when "00100000011100",
                      106 when "00100000011101",
                      106 when "00100000011110",
                      106 when "00100000011111",
                      106 when "00100000100000",
                      106 when "00100000100001",
                      106 when "00100000100010",
                      105 when "00100000100011",
                      105 when "00100000100100",
                      105 when "00100000100101",
                      105 when "00100000100110",
                      105 when "00100000100111",
                      105 when "00100000101000",
                      105 when "00100000101001",
                      105 when "00100000101010",
                      105 when "00100000101011",
                      105 when "00100000101100",
                      105 when "00100000101101",
                      105 when "00100000101110",
                      105 when "00100000101111",
                      105 when "00100000110000",
                      105 when "00100000110001",
                      105 when "00100000110010",
                      105 when "00100000110011",
                      105 when "00100000110100",
                      105 when "00100000110101",
                      105 when "00100000110110",
                      104 when "00100000110111",
                      104 when "00100000111000",
                      104 when "00100000111001",
                      104 when "00100000111010",
                      104 when "00100000111011",
                      104 when "00100000111100",
                      104 when "00100000111101",
                      104 when "00100000111110",
                      104 when "00100000111111",
                      104 when "00100001000000",
                      104 when "00100001000001",
                      104 when "00100001000010",
                      104 when "00100001000011",
                      104 when "00100001000100",
                      104 when "00100001000101",
                      104 when "00100001000110",
                      104 when "00100001000111",
                      104 when "00100001001000",
                      104 when "00100001001001",
                      104 when "00100001001010",
                      103 when "00100001001011",
                      103 when "00100001001100",
                      103 when "00100001001101",
                      103 when "00100001001110",
                      103 when "00100001001111",
                      103 when "00100001010000",
                      103 when "00100001010001",
                      103 when "00100001010010",
                      103 when "00100001010011",
                      103 when "00100001010100",
                      103 when "00100001010101",
                      103 when "00100001010110",
                      103 when "00100001010111",
                      103 when "00100001011000",
                      103 when "00100001011001",
                      103 when "00100001011010",
                      103 when "00100001011011",
                      103 when "00100001011100",
                      103 when "00100001011101",
                      103 when "00100001011110",
                      103 when "00100001011111",
                      102 when "00100001100000",
                      102 when "00100001100001",
                      102 when "00100001100010",
                      102 when "00100001100011",
                      102 when "00100001100100",
                      102 when "00100001100101",
                      102 when "00100001100110",
                      102 when "00100001100111",
                      102 when "00100001101000",
                      102 when "00100001101001",
                      102 when "00100001101010",
                      102 when "00100001101011",
                      102 when "00100001101100",
                      102 when "00100001101101",
                      102 when "00100001101110",
                      102 when "00100001101111",
                      102 when "00100001110000",
                      102 when "00100001110001",
                      102 when "00100001110010",
                      102 when "00100001110011",
                      102 when "00100001110100",
                      101 when "00100001110101",
                      101 when "00100001110110",
                      101 when "00100001110111",
                      101 when "00100001111000",
                      101 when "00100001111001",
                      101 when "00100001111010",
                      101 when "00100001111011",
                      101 when "00100001111100",
                      101 when "00100001111101",
                      101 when "00100001111110",
                      101 when "00100001111111",
                      101 when "00100010000000",
                      101 when "00100010000001",
                      101 when "00100010000010",
                      101 when "00100010000011",
                      101 when "00100010000100",
                      101 when "00100010000101",
                      101 when "00100010000110",
                      101 when "00100010000111",
                      101 when "00100010001000",
                      101 when "00100010001001",
                      101 when "00100010001010",
                      100 when "00100010001011",
                      100 when "00100010001100",
                      100 when "00100010001101",
                      100 when "00100010001110",
                      100 when "00100010001111",
                      100 when "00100010010000",
                      100 when "00100010010001",
                      100 when "00100010010010",
                      100 when "00100010010011",
                      100 when "00100010010100",
                      100 when "00100010010101",
                      100 when "00100010010110",
                      100 when "00100010010111",
                      100 when "00100010011000",
                      100 when "00100010011001",
                      100 when "00100010011010",
                      100 when "00100010011011",
                      100 when "00100010011100",
                      100 when "00100010011101",
                      100 when "00100010011110",
                      100 when "00100010011111",
                      100 when "00100010100000",
                      99 when "00100010100001",
                      99 when "00100010100010",
                      99 when "00100010100011",
                      99 when "00100010100100",
                      99 when "00100010100101",
                      99 when "00100010100110",
                      99 when "00100010100111",
                      99 when "00100010101000",
                      99 when "00100010101001",
                      99 when "00100010101010",
                      99 when "00100010101011",
                      99 when "00100010101100",
                      99 when "00100010101101",
                      99 when "00100010101110",
                      99 when "00100010101111",
                      99 when "00100010110000",
                      99 when "00100010110001",
                      99 when "00100010110010",
                      99 when "00100010110011",
                      99 when "00100010110100",
                      99 when "00100010110101",
                      99 when "00100010110110",
                      98 when "00100010110111",
                      98 when "00100010111000",
                      98 when "00100010111001",
                      98 when "00100010111010",
                      98 when "00100010111011",
                      98 when "00100010111100",
                      98 when "00100010111101",
                      98 when "00100010111110",
                      98 when "00100010111111",
                      98 when "00100011000000",
                      98 when "00100011000001",
                      98 when "00100011000010",
                      98 when "00100011000011",
                      98 when "00100011000100",
                      98 when "00100011000101",
                      98 when "00100011000110",
                      98 when "00100011000111",
                      98 when "00100011001000",
                      98 when "00100011001001",
                      98 when "00100011001010",
                      98 when "00100011001011",
                      98 when "00100011001100",
                      98 when "00100011001101",
                      97 when "00100011001110",
                      97 when "00100011001111",
                      97 when "00100011010000",
                      97 when "00100011010001",
                      97 when "00100011010010",
                      97 when "00100011010011",
                      97 when "00100011010100",
                      97 when "00100011010101",
                      97 when "00100011010110",
                      97 when "00100011010111",
                      97 when "00100011011000",
                      97 when "00100011011001",
                      97 when "00100011011010",
                      97 when "00100011011011",
                      97 when "00100011011100",
                      97 when "00100011011101",
                      97 when "00100011011110",
                      97 when "00100011011111",
                      97 when "00100011100000",
                      97 when "00100011100001",
                      97 when "00100011100010",
                      97 when "00100011100011",
                      97 when "00100011100100",
                      96 when "00100011100101",
                      96 when "00100011100110",
                      96 when "00100011100111",
                      96 when "00100011101000",
                      96 when "00100011101001",
                      96 when "00100011101010",
                      96 when "00100011101011",
                      96 when "00100011101100",
                      96 when "00100011101101",
                      96 when "00100011101110",
                      96 when "00100011101111",
                      96 when "00100011110000",
                      96 when "00100011110001",
                      96 when "00100011110010",
                      96 when "00100011110011",
                      96 when "00100011110100",
                      96 when "00100011110101",
                      96 when "00100011110110",
                      96 when "00100011110111",
                      96 when "00100011111000",
                      96 when "00100011111001",
                      96 when "00100011111010",
                      96 when "00100011111011",
                      96 when "00100011111100",
                      95 when "00100011111101",
                      95 when "00100011111110",
                      95 when "00100011111111",
                      95 when "00100100000000",
                      95 when "00100100000001",
                      95 when "00100100000010",
                      95 when "00100100000011",
                      95 when "00100100000100",
                      95 when "00100100000101",
                      95 when "00100100000110",
                      95 when "00100100000111",
                      95 when "00100100001000",
                      95 when "00100100001001",
                      95 when "00100100001010",
                      95 when "00100100001011",
                      95 when "00100100001100",
                      95 when "00100100001101",
                      95 when "00100100001110",
                      95 when "00100100001111",
                      95 when "00100100010000",
                      95 when "00100100010001",
                      95 when "00100100010010",
                      95 when "00100100010011",
                      95 when "00100100010100",
                      95 when "00100100010101",
                      94 when "00100100010110",
                      94 when "00100100010111",
                      94 when "00100100011000",
                      94 when "00100100011001",
                      94 when "00100100011010",
                      94 when "00100100011011",
                      94 when "00100100011100",
                      94 when "00100100011101",
                      94 when "00100100011110",
                      94 when "00100100011111",
                      94 when "00100100100000",
                      94 when "00100100100001",
                      94 when "00100100100010",
                      94 when "00100100100011",
                      94 when "00100100100100",
                      94 when "00100100100101",
                      94 when "00100100100110",
                      94 when "00100100100111",
                      94 when "00100100101000",
                      94 when "00100100101001",
                      94 when "00100100101010",
                      94 when "00100100101011",
                      94 when "00100100101100",
                      94 when "00100100101101",
                      94 when "00100100101110",
                      93 when "00100100101111",
                      93 when "00100100110000",
                      93 when "00100100110001",
                      93 when "00100100110010",
                      93 when "00100100110011",
                      93 when "00100100110100",
                      93 when "00100100110101",
                      93 when "00100100110110",
                      93 when "00100100110111",
                      93 when "00100100111000",
                      93 when "00100100111001",
                      93 when "00100100111010",
                      93 when "00100100111011",
                      93 when "00100100111100",
                      93 when "00100100111101",
                      93 when "00100100111110",
                      93 when "00100100111111",
                      93 when "00100101000000",
                      93 when "00100101000001",
                      93 when "00100101000010",
                      93 when "00100101000011",
                      93 when "00100101000100",
                      93 when "00100101000101",
                      93 when "00100101000110",
                      93 when "00100101000111",
                      92 when "00100101001000",
                      92 when "00100101001001",
                      92 when "00100101001010",
                      92 when "00100101001011",
                      92 when "00100101001100",
                      92 when "00100101001101",
                      92 when "00100101001110",
                      92 when "00100101001111",
                      92 when "00100101010000",
                      92 when "00100101010001",
                      92 when "00100101010010",
                      92 when "00100101010011",
                      92 when "00100101010100",
                      92 when "00100101010101",
                      92 when "00100101010110",
                      92 when "00100101010111",
                      92 when "00100101011000",
                      92 when "00100101011001",
                      92 when "00100101011010",
                      92 when "00100101011011",
                      92 when "00100101011100",
                      92 when "00100101011101",
                      92 when "00100101011110",
                      92 when "00100101011111",
                      92 when "00100101100000",
                      92 when "00100101100001",
                      91 when "00100101100010",
                      91 when "00100101100011",
                      91 when "00100101100100",
                      91 when "00100101100101",
                      91 when "00100101100110",
                      91 when "00100101100111",
                      91 when "00100101101000",
                      91 when "00100101101001",
                      91 when "00100101101010",
                      91 when "00100101101011",
                      91 when "00100101101100",
                      91 when "00100101101101",
                      91 when "00100101101110",
                      91 when "00100101101111",
                      91 when "00100101110000",
                      91 when "00100101110001",
                      91 when "00100101110010",
                      91 when "00100101110011",
                      91 when "00100101110100",
                      91 when "00100101110101",
                      91 when "00100101110110",
                      91 when "00100101110111",
                      91 when "00100101111000",
                      91 when "00100101111001",
                      91 when "00100101111010",
                      91 when "00100101111011",
                      90 when "00100101111100",
                      90 when "00100101111101",
                      90 when "00100101111110",
                      90 when "00100101111111",
                      90 when "00100110000000",
                      90 when "00100110000001",
                      90 when "00100110000010",
                      90 when "00100110000011",
                      90 when "00100110000100",
                      90 when "00100110000101",
                      90 when "00100110000110",
                      90 when "00100110000111",
                      90 when "00100110001000",
                      90 when "00100110001001",
                      90 when "00100110001010",
                      90 when "00100110001011",
                      90 when "00100110001100",
                      90 when "00100110001101",
                      90 when "00100110001110",
                      90 when "00100110001111",
                      90 when "00100110010000",
                      90 when "00100110010001",
                      90 when "00100110010010",
                      90 when "00100110010011",
                      90 when "00100110010100",
                      90 when "00100110010101",
                      90 when "00100110010110",
                      90 when "00100110010111",
                      89 when "00100110011000",
                      89 when "00100110011001",
                      89 when "00100110011010",
                      89 when "00100110011011",
                      89 when "00100110011100",
                      89 when "00100110011101",
                      89 when "00100110011110",
                      89 when "00100110011111",
                      89 when "00100110100000",
                      89 when "00100110100001",
                      89 when "00100110100010",
                      89 when "00100110100011",
                      89 when "00100110100100",
                      89 when "00100110100101",
                      89 when "00100110100110",
                      89 when "00100110100111",
                      89 when "00100110101000",
                      89 when "00100110101001",
                      89 when "00100110101010",
                      89 when "00100110101011",
                      89 when "00100110101100",
                      89 when "00100110101101",
                      89 when "00100110101110",
                      89 when "00100110101111",
                      89 when "00100110110000",
                      89 when "00100110110001",
                      89 when "00100110110010",
                      88 when "00100110110011",
                      88 when "00100110110100",
                      88 when "00100110110101",
                      88 when "00100110110110",
                      88 when "00100110110111",
                      88 when "00100110111000",
                      88 when "00100110111001",
                      88 when "00100110111010",
                      88 when "00100110111011",
                      88 when "00100110111100",
                      88 when "00100110111101",
                      88 when "00100110111110",
                      88 when "00100110111111",
                      88 when "00100111000000",
                      88 when "00100111000001",
                      88 when "00100111000010",
                      88 when "00100111000011",
                      88 when "00100111000100",
                      88 when "00100111000101",
                      88 when "00100111000110",
                      88 when "00100111000111",
                      88 when "00100111001000",
                      88 when "00100111001001",
                      88 when "00100111001010",
                      88 when "00100111001011",
                      88 when "00100111001100",
                      88 when "00100111001101",
                      88 when "00100111001110",
                      88 when "00100111001111",
                      87 when "00100111010000",
                      87 when "00100111010001",
                      87 when "00100111010010",
                      87 when "00100111010011",
                      87 when "00100111010100",
                      87 when "00100111010101",
                      87 when "00100111010110",
                      87 when "00100111010111",
                      87 when "00100111011000",
                      87 when "00100111011001",
                      87 when "00100111011010",
                      87 when "00100111011011",
                      87 when "00100111011100",
                      87 when "00100111011101",
                      87 when "00100111011110",
                      87 when "00100111011111",
                      87 when "00100111100000",
                      87 when "00100111100001",
                      87 when "00100111100010",
                      87 when "00100111100011",
                      87 when "00100111100100",
                      87 when "00100111100101",
                      87 when "00100111100110",
                      87 when "00100111100111",
                      87 when "00100111101000",
                      87 when "00100111101001",
                      87 when "00100111101010",
                      87 when "00100111101011",
                      87 when "00100111101100",
                      86 when "00100111101101",
                      86 when "00100111101110",
                      86 when "00100111101111",
                      86 when "00100111110000",
                      86 when "00100111110001",
                      86 when "00100111110010",
                      86 when "00100111110011",
                      86 when "00100111110100",
                      86 when "00100111110101",
                      86 when "00100111110110",
                      86 when "00100111110111",
                      86 when "00100111111000",
                      86 when "00100111111001",
                      86 when "00100111111010",
                      86 when "00100111111011",
                      86 when "00100111111100",
                      86 when "00100111111101",
                      86 when "00100111111110",
                      86 when "00100111111111",
                      86 when "00101000000000",
                      86 when "00101000000001",
                      86 when "00101000000010",
                      86 when "00101000000011",
                      86 when "00101000000100",
                      86 when "00101000000101",
                      86 when "00101000000110",
                      86 when "00101000000111",
                      86 when "00101000001000",
                      86 when "00101000001001",
                      85 when "00101000001010",
                      85 when "00101000001011",
                      85 when "00101000001100",
                      85 when "00101000001101",
                      85 when "00101000001110",
                      85 when "00101000001111",
                      85 when "00101000010000",
                      85 when "00101000010001",
                      85 when "00101000010010",
                      85 when "00101000010011",
                      85 when "00101000010100",
                      85 when "00101000010101",
                      85 when "00101000010110",
                      85 when "00101000010111",
                      85 when "00101000011000",
                      85 when "00101000011001",
                      85 when "00101000011010",
                      85 when "00101000011011",
                      85 when "00101000011100",
                      85 when "00101000011101",
                      85 when "00101000011110",
                      85 when "00101000011111",
                      85 when "00101000100000",
                      85 when "00101000100001",
                      85 when "00101000100010",
                      85 when "00101000100011",
                      85 when "00101000100100",
                      85 when "00101000100101",
                      85 when "00101000100110",
                      85 when "00101000100111",
                      85 when "00101000101000",
                      84 when "00101000101001",
                      84 when "00101000101010",
                      84 when "00101000101011",
                      84 when "00101000101100",
                      84 when "00101000101101",
                      84 when "00101000101110",
                      84 when "00101000101111",
                      84 when "00101000110000",
                      84 when "00101000110001",
                      84 when "00101000110010",
                      84 when "00101000110011",
                      84 when "00101000110100",
                      84 when "00101000110101",
                      84 when "00101000110110",
                      84 when "00101000110111",
                      84 when "00101000111000",
                      84 when "00101000111001",
                      84 when "00101000111010",
                      84 when "00101000111011",
                      84 when "00101000111100",
                      84 when "00101000111101",
                      84 when "00101000111110",
                      84 when "00101000111111",
                      84 when "00101001000000",
                      84 when "00101001000001",
                      84 when "00101001000010",
                      84 when "00101001000011",
                      84 when "00101001000100",
                      84 when "00101001000101",
                      84 when "00101001000110",
                      84 when "00101001000111",
                      83 when "00101001001000",
                      83 when "00101001001001",
                      83 when "00101001001010",
                      83 when "00101001001011",
                      83 when "00101001001100",
                      83 when "00101001001101",
                      83 when "00101001001110",
                      83 when "00101001001111",
                      83 when "00101001010000",
                      83 when "00101001010001",
                      83 when "00101001010010",
                      83 when "00101001010011",
                      83 when "00101001010100",
                      83 when "00101001010101",
                      83 when "00101001010110",
                      83 when "00101001010111",
                      83 when "00101001011000",
                      83 when "00101001011001",
                      83 when "00101001011010",
                      83 when "00101001011011",
                      83 when "00101001011100",
                      83 when "00101001011101",
                      83 when "00101001011110",
                      83 when "00101001011111",
                      83 when "00101001100000",
                      83 when "00101001100001",
                      83 when "00101001100010",
                      83 when "00101001100011",
                      83 when "00101001100100",
                      83 when "00101001100101",
                      83 when "00101001100110",
                      83 when "00101001100111",
                      82 when "00101001101000",
                      82 when "00101001101001",
                      82 when "00101001101010",
                      82 when "00101001101011",
                      82 when "00101001101100",
                      82 when "00101001101101",
                      82 when "00101001101110",
                      82 when "00101001101111",
                      82 when "00101001110000",
                      82 when "00101001110001",
                      82 when "00101001110010",
                      82 when "00101001110011",
                      82 when "00101001110100",
                      82 when "00101001110101",
                      82 when "00101001110110",
                      82 when "00101001110111",
                      82 when "00101001111000",
                      82 when "00101001111001",
                      82 when "00101001111010",
                      82 when "00101001111011",
                      82 when "00101001111100",
                      82 when "00101001111101",
                      82 when "00101001111110",
                      82 when "00101001111111",
                      82 when "00101010000000",
                      82 when "00101010000001",
                      82 when "00101010000010",
                      82 when "00101010000011",
                      82 when "00101010000100",
                      82 when "00101010000101",
                      82 when "00101010000110",
                      82 when "00101010000111",
                      82 when "00101010001000",
                      81 when "00101010001001",
                      81 when "00101010001010",
                      81 when "00101010001011",
                      81 when "00101010001100",
                      81 when "00101010001101",
                      81 when "00101010001110",
                      81 when "00101010001111",
                      81 when "00101010010000",
                      81 when "00101010010001",
                      81 when "00101010010010",
                      81 when "00101010010011",
                      81 when "00101010010100",
                      81 when "00101010010101",
                      81 when "00101010010110",
                      81 when "00101010010111",
                      81 when "00101010011000",
                      81 when "00101010011001",
                      81 when "00101010011010",
                      81 when "00101010011011",
                      81 when "00101010011100",
                      81 when "00101010011101",
                      81 when "00101010011110",
                      81 when "00101010011111",
                      81 when "00101010100000",
                      81 when "00101010100001",
                      81 when "00101010100010",
                      81 when "00101010100011",
                      81 when "00101010100100",
                      81 when "00101010100101",
                      81 when "00101010100110",
                      81 when "00101010100111",
                      81 when "00101010101000",
                      81 when "00101010101001",
                      80 when "00101010101010",
                      80 when "00101010101011",
                      80 when "00101010101100",
                      80 when "00101010101101",
                      80 when "00101010101110",
                      80 when "00101010101111",
                      80 when "00101010110000",
                      80 when "00101010110001",
                      80 when "00101010110010",
                      80 when "00101010110011",
                      80 when "00101010110100",
                      80 when "00101010110101",
                      80 when "00101010110110",
                      80 when "00101010110111",
                      80 when "00101010111000",
                      80 when "00101010111001",
                      80 when "00101010111010",
                      80 when "00101010111011",
                      80 when "00101010111100",
                      80 when "00101010111101",
                      80 when "00101010111110",
                      80 when "00101010111111",
                      80 when "00101011000000",
                      80 when "00101011000001",
                      80 when "00101011000010",
                      80 when "00101011000011",
                      80 when "00101011000100",
                      80 when "00101011000101",
                      80 when "00101011000110",
                      80 when "00101011000111",
                      80 when "00101011001000",
                      80 when "00101011001001",
                      80 when "00101011001010",
                      80 when "00101011001011",
                      79 when "00101011001100",
                      79 when "00101011001101",
                      79 when "00101011001110",
                      79 when "00101011001111",
                      79 when "00101011010000",
                      79 when "00101011010001",
                      79 when "00101011010010",
                      79 when "00101011010011",
                      79 when "00101011010100",
                      79 when "00101011010101",
                      79 when "00101011010110",
                      79 when "00101011010111",
                      79 when "00101011011000",
                      79 when "00101011011001",
                      79 when "00101011011010",
                      79 when "00101011011011",
                      79 when "00101011011100",
                      79 when "00101011011101",
                      79 when "00101011011110",
                      79 when "00101011011111",
                      79 when "00101011100000",
                      79 when "00101011100001",
                      79 when "00101011100010",
                      79 when "00101011100011",
                      79 when "00101011100100",
                      79 when "00101011100101",
                      79 when "00101011100110",
                      79 when "00101011100111",
                      79 when "00101011101000",
                      79 when "00101011101001",
                      79 when "00101011101010",
                      79 when "00101011101011",
                      79 when "00101011101100",
                      79 when "00101011101101",
                      79 when "00101011101110",
                      79 when "00101011101111",
                      78 when "00101011110000",
                      78 when "00101011110001",
                      78 when "00101011110010",
                      78 when "00101011110011",
                      78 when "00101011110100",
                      78 when "00101011110101",
                      78 when "00101011110110",
                      78 when "00101011110111",
                      78 when "00101011111000",
                      78 when "00101011111001",
                      78 when "00101011111010",
                      78 when "00101011111011",
                      78 when "00101011111100",
                      78 when "00101011111101",
                      78 when "00101011111110",
                      78 when "00101011111111",
                      78 when "00101100000000",
                      78 when "00101100000001",
                      78 when "00101100000010",
                      78 when "00101100000011",
                      78 when "00101100000100",
                      78 when "00101100000101",
                      78 when "00101100000110",
                      78 when "00101100000111",
                      78 when "00101100001000",
                      78 when "00101100001001",
                      78 when "00101100001010",
                      78 when "00101100001011",
                      78 when "00101100001100",
                      78 when "00101100001101",
                      78 when "00101100001110",
                      78 when "00101100001111",
                      78 when "00101100010000",
                      78 when "00101100010001",
                      78 when "00101100010010",
                      78 when "00101100010011",
                      77 when "00101100010100",
                      77 when "00101100010101",
                      77 when "00101100010110",
                      77 when "00101100010111",
                      77 when "00101100011000",
                      77 when "00101100011001",
                      77 when "00101100011010",
                      77 when "00101100011011",
                      77 when "00101100011100",
                      77 when "00101100011101",
                      77 when "00101100011110",
                      77 when "00101100011111",
                      77 when "00101100100000",
                      77 when "00101100100001",
                      77 when "00101100100010",
                      77 when "00101100100011",
                      77 when "00101100100100",
                      77 when "00101100100101",
                      77 when "00101100100110",
                      77 when "00101100100111",
                      77 when "00101100101000",
                      77 when "00101100101001",
                      77 when "00101100101010",
                      77 when "00101100101011",
                      77 when "00101100101100",
                      77 when "00101100101101",
                      77 when "00101100101110",
                      77 when "00101100101111",
                      77 when "00101100110000",
                      77 when "00101100110001",
                      77 when "00101100110010",
                      77 when "00101100110011",
                      77 when "00101100110100",
                      77 when "00101100110101",
                      77 when "00101100110110",
                      77 when "00101100110111",
                      77 when "00101100111000",
                      76 when "00101100111001",
                      76 when "00101100111010",
                      76 when "00101100111011",
                      76 when "00101100111100",
                      76 when "00101100111101",
                      76 when "00101100111110",
                      76 when "00101100111111",
                      76 when "00101101000000",
                      76 when "00101101000001",
                      76 when "00101101000010",
                      76 when "00101101000011",
                      76 when "00101101000100",
                      76 when "00101101000101",
                      76 when "00101101000110",
                      76 when "00101101000111",
                      76 when "00101101001000",
                      76 when "00101101001001",
                      76 when "00101101001010",
                      76 when "00101101001011",
                      76 when "00101101001100",
                      76 when "00101101001101",
                      76 when "00101101001110",
                      76 when "00101101001111",
                      76 when "00101101010000",
                      76 when "00101101010001",
                      76 when "00101101010010",
                      76 when "00101101010011",
                      76 when "00101101010100",
                      76 when "00101101010101",
                      76 when "00101101010110",
                      76 when "00101101010111",
                      76 when "00101101011000",
                      76 when "00101101011001",
                      76 when "00101101011010",
                      76 when "00101101011011",
                      76 when "00101101011100",
                      76 when "00101101011101",
                      76 when "00101101011110",
                      75 when "00101101011111",
                      75 when "00101101100000",
                      75 when "00101101100001",
                      75 when "00101101100010",
                      75 when "00101101100011",
                      75 when "00101101100100",
                      75 when "00101101100101",
                      75 when "00101101100110",
                      75 when "00101101100111",
                      75 when "00101101101000",
                      75 when "00101101101001",
                      75 when "00101101101010",
                      75 when "00101101101011",
                      75 when "00101101101100",
                      75 when "00101101101101",
                      75 when "00101101101110",
                      75 when "00101101101111",
                      75 when "00101101110000",
                      75 when "00101101110001",
                      75 when "00101101110010",
                      75 when "00101101110011",
                      75 when "00101101110100",
                      75 when "00101101110101",
                      75 when "00101101110110",
                      75 when "00101101110111",
                      75 when "00101101111000",
                      75 when "00101101111001",
                      75 when "00101101111010",
                      75 when "00101101111011",
                      75 when "00101101111100",
                      75 when "00101101111101",
                      75 when "00101101111110",
                      75 when "00101101111111",
                      75 when "00101110000000",
                      75 when "00101110000001",
                      75 when "00101110000010",
                      75 when "00101110000011",
                      75 when "00101110000100",
                      75 when "00101110000101",
                      74 when "00101110000110",
                      74 when "00101110000111",
                      74 when "00101110001000",
                      74 when "00101110001001",
                      74 when "00101110001010",
                      74 when "00101110001011",
                      74 when "00101110001100",
                      74 when "00101110001101",
                      74 when "00101110001110",
                      74 when "00101110001111",
                      74 when "00101110010000",
                      74 when "00101110010001",
                      74 when "00101110010010",
                      74 when "00101110010011",
                      74 when "00101110010100",
                      74 when "00101110010101",
                      74 when "00101110010110",
                      74 when "00101110010111",
                      74 when "00101110011000",
                      74 when "00101110011001",
                      74 when "00101110011010",
                      74 when "00101110011011",
                      74 when "00101110011100",
                      74 when "00101110011101",
                      74 when "00101110011110",
                      74 when "00101110011111",
                      74 when "00101110100000",
                      74 when "00101110100001",
                      74 when "00101110100010",
                      74 when "00101110100011",
                      74 when "00101110100100",
                      74 when "00101110100101",
                      74 when "00101110100110",
                      74 when "00101110100111",
                      74 when "00101110101000",
                      74 when "00101110101001",
                      74 when "00101110101010",
                      74 when "00101110101011",
                      74 when "00101110101100",
                      74 when "00101110101101",
                      73 when "00101110101110",
                      73 when "00101110101111",
                      73 when "00101110110000",
                      73 when "00101110110001",
                      73 when "00101110110010",
                      73 when "00101110110011",
                      73 when "00101110110100",
                      73 when "00101110110101",
                      73 when "00101110110110",
                      73 when "00101110110111",
                      73 when "00101110111000",
                      73 when "00101110111001",
                      73 when "00101110111010",
                      73 when "00101110111011",
                      73 when "00101110111100",
                      73 when "00101110111101",
                      73 when "00101110111110",
                      73 when "00101110111111",
                      73 when "00101111000000",
                      73 when "00101111000001",
                      73 when "00101111000010",
                      73 when "00101111000011",
                      73 when "00101111000100",
                      73 when "00101111000101",
                      73 when "00101111000110",
                      73 when "00101111000111",
                      73 when "00101111001000",
                      73 when "00101111001001",
                      73 when "00101111001010",
                      73 when "00101111001011",
                      73 when "00101111001100",
                      73 when "00101111001101",
                      73 when "00101111001110",
                      73 when "00101111001111",
                      73 when "00101111010000",
                      73 when "00101111010001",
                      73 when "00101111010010",
                      73 when "00101111010011",
                      73 when "00101111010100",
                      73 when "00101111010101",
                      73 when "00101111010110",
                      72 when "00101111010111",
                      72 when "00101111011000",
                      72 when "00101111011001",
                      72 when "00101111011010",
                      72 when "00101111011011",
                      72 when "00101111011100",
                      72 when "00101111011101",
                      72 when "00101111011110",
                      72 when "00101111011111",
                      72 when "00101111100000",
                      72 when "00101111100001",
                      72 when "00101111100010",
                      72 when "00101111100011",
                      72 when "00101111100100",
                      72 when "00101111100101",
                      72 when "00101111100110",
                      72 when "00101111100111",
                      72 when "00101111101000",
                      72 when "00101111101001",
                      72 when "00101111101010",
                      72 when "00101111101011",
                      72 when "00101111101100",
                      72 when "00101111101101",
                      72 when "00101111101110",
                      72 when "00101111101111",
                      72 when "00101111110000",
                      72 when "00101111110001",
                      72 when "00101111110010",
                      72 when "00101111110011",
                      72 when "00101111110100",
                      72 when "00101111110101",
                      72 when "00101111110110",
                      72 when "00101111110111",
                      72 when "00101111111000",
                      72 when "00101111111001",
                      72 when "00101111111010",
                      72 when "00101111111011",
                      72 when "00101111111100",
                      72 when "00101111111101",
                      72 when "00101111111110",
                      72 when "00101111111111",
                      72 when "00110000000000",
                      72 when "00110000000001",
                      71 when "00110000000010",
                      71 when "00110000000011",
                      71 when "00110000000100",
                      71 when "00110000000101",
                      71 when "00110000000110",
                      71 when "00110000000111",
                      71 when "00110000001000",
                      71 when "00110000001001",
                      71 when "00110000001010",
                      71 when "00110000001011",
                      71 when "00110000001100",
                      71 when "00110000001101",
                      71 when "00110000001110",
                      71 when "00110000001111",
                      71 when "00110000010000",
                      71 when "00110000010001",
                      71 when "00110000010010",
                      71 when "00110000010011",
                      71 when "00110000010100",
                      71 when "00110000010101",
                      71 when "00110000010110",
                      71 when "00110000010111",
                      71 when "00110000011000",
                      71 when "00110000011001",
                      71 when "00110000011010",
                      71 when "00110000011011",
                      71 when "00110000011100",
                      71 when "00110000011101",
                      71 when "00110000011110",
                      71 when "00110000011111",
                      71 when "00110000100000",
                      71 when "00110000100001",
                      71 when "00110000100010",
                      71 when "00110000100011",
                      71 when "00110000100100",
                      71 when "00110000100101",
                      71 when "00110000100110",
                      71 when "00110000100111",
                      71 when "00110000101000",
                      71 when "00110000101001",
                      71 when "00110000101010",
                      71 when "00110000101011",
                      71 when "00110000101100",
                      70 when "00110000101101",
                      70 when "00110000101110",
                      70 when "00110000101111",
                      70 when "00110000110000",
                      70 when "00110000110001",
                      70 when "00110000110010",
                      70 when "00110000110011",
                      70 when "00110000110100",
                      70 when "00110000110101",
                      70 when "00110000110110",
                      70 when "00110000110111",
                      70 when "00110000111000",
                      70 when "00110000111001",
                      70 when "00110000111010",
                      70 when "00110000111011",
                      70 when "00110000111100",
                      70 when "00110000111101",
                      70 when "00110000111110",
                      70 when "00110000111111",
                      70 when "00110001000000",
                      70 when "00110001000001",
                      70 when "00110001000010",
                      70 when "00110001000011",
                      70 when "00110001000100",
                      70 when "00110001000101",
                      70 when "00110001000110",
                      70 when "00110001000111",
                      70 when "00110001001000",
                      70 when "00110001001001",
                      70 when "00110001001010",
                      70 when "00110001001011",
                      70 when "00110001001100",
                      70 when "00110001001101",
                      70 when "00110001001110",
                      70 when "00110001001111",
                      70 when "00110001010000",
                      70 when "00110001010001",
                      70 when "00110001010010",
                      70 when "00110001010011",
                      70 when "00110001010100",
                      70 when "00110001010101",
                      70 when "00110001010110",
                      70 when "00110001010111",
                      70 when "00110001011000",
                      70 when "00110001011001",
                      69 when "00110001011010",
                      69 when "00110001011011",
                      69 when "00110001011100",
                      69 when "00110001011101",
                      69 when "00110001011110",
                      69 when "00110001011111",
                      69 when "00110001100000",
                      69 when "00110001100001",
                      69 when "00110001100010",
                      69 when "00110001100011",
                      69 when "00110001100100",
                      69 when "00110001100101",
                      69 when "00110001100110",
                      69 when "00110001100111",
                      69 when "00110001101000",
                      69 when "00110001101001",
                      69 when "00110001101010",
                      69 when "00110001101011",
                      69 when "00110001101100",
                      69 when "00110001101101",
                      69 when "00110001101110",
                      69 when "00110001101111",
                      69 when "00110001110000",
                      69 when "00110001110001",
                      69 when "00110001110010",
                      69 when "00110001110011",
                      69 when "00110001110100",
                      69 when "00110001110101",
                      69 when "00110001110110",
                      69 when "00110001110111",
                      69 when "00110001111000",
                      69 when "00110001111001",
                      69 when "00110001111010",
                      69 when "00110001111011",
                      69 when "00110001111100",
                      69 when "00110001111101",
                      69 when "00110001111110",
                      69 when "00110001111111",
                      69 when "00110010000000",
                      69 when "00110010000001",
                      69 when "00110010000010",
                      69 when "00110010000011",
                      69 when "00110010000100",
                      69 when "00110010000101",
                      69 when "00110010000110",
                      69 when "00110010000111",
                      68 when "00110010001000",
                      68 when "00110010001001",
                      68 when "00110010001010",
                      68 when "00110010001011",
                      68 when "00110010001100",
                      68 when "00110010001101",
                      68 when "00110010001110",
                      68 when "00110010001111",
                      68 when "00110010010000",
                      68 when "00110010010001",
                      68 when "00110010010010",
                      68 when "00110010010011",
                      68 when "00110010010100",
                      68 when "00110010010101",
                      68 when "00110010010110",
                      68 when "00110010010111",
                      68 when "00110010011000",
                      68 when "00110010011001",
                      68 when "00110010011010",
                      68 when "00110010011011",
                      68 when "00110010011100",
                      68 when "00110010011101",
                      68 when "00110010011110",
                      68 when "00110010011111",
                      68 when "00110010100000",
                      68 when "00110010100001",
                      68 when "00110010100010",
                      68 when "00110010100011",
                      68 when "00110010100100",
                      68 when "00110010100101",
                      68 when "00110010100110",
                      68 when "00110010100111",
                      68 when "00110010101000",
                      68 when "00110010101001",
                      68 when "00110010101010",
                      68 when "00110010101011",
                      68 when "00110010101100",
                      68 when "00110010101101",
                      68 when "00110010101110",
                      68 when "00110010101111",
                      68 when "00110010110000",
                      68 when "00110010110001",
                      68 when "00110010110010",
                      68 when "00110010110011",
                      68 when "00110010110100",
                      68 when "00110010110101",
                      68 when "00110010110110",
                      68 when "00110010110111",
                      67 when "00110010111000",
                      67 when "00110010111001",
                      67 when "00110010111010",
                      67 when "00110010111011",
                      67 when "00110010111100",
                      67 when "00110010111101",
                      67 when "00110010111110",
                      67 when "00110010111111",
                      67 when "00110011000000",
                      67 when "00110011000001",
                      67 when "00110011000010",
                      67 when "00110011000011",
                      67 when "00110011000100",
                      67 when "00110011000101",
                      67 when "00110011000110",
                      67 when "00110011000111",
                      67 when "00110011001000",
                      67 when "00110011001001",
                      67 when "00110011001010",
                      67 when "00110011001011",
                      67 when "00110011001100",
                      67 when "00110011001101",
                      67 when "00110011001110",
                      67 when "00110011001111",
                      67 when "00110011010000",
                      67 when "00110011010001",
                      67 when "00110011010010",
                      67 when "00110011010011",
                      67 when "00110011010100",
                      67 when "00110011010101",
                      67 when "00110011010110",
                      67 when "00110011010111",
                      67 when "00110011011000",
                      67 when "00110011011001",
                      67 when "00110011011010",
                      67 when "00110011011011",
                      67 when "00110011011100",
                      67 when "00110011011101",
                      67 when "00110011011110",
                      67 when "00110011011111",
                      67 when "00110011100000",
                      67 when "00110011100001",
                      67 when "00110011100010",
                      67 when "00110011100011",
                      67 when "00110011100100",
                      67 when "00110011100101",
                      67 when "00110011100110",
                      67 when "00110011100111",
                      67 when "00110011101000",
                      66 when "00110011101001",
                      66 when "00110011101010",
                      66 when "00110011101011",
                      66 when "00110011101100",
                      66 when "00110011101101",
                      66 when "00110011101110",
                      66 when "00110011101111",
                      66 when "00110011110000",
                      66 when "00110011110001",
                      66 when "00110011110010",
                      66 when "00110011110011",
                      66 when "00110011110100",
                      66 when "00110011110101",
                      66 when "00110011110110",
                      66 when "00110011110111",
                      66 when "00110011111000",
                      66 when "00110011111001",
                      66 when "00110011111010",
                      66 when "00110011111011",
                      66 when "00110011111100",
                      66 when "00110011111101",
                      66 when "00110011111110",
                      66 when "00110011111111",
                      66 when "00110100000000",
                      66 when "00110100000001",
                      66 when "00110100000010",
                      66 when "00110100000011",
                      66 when "00110100000100",
                      66 when "00110100000101",
                      66 when "00110100000110",
                      66 when "00110100000111",
                      66 when "00110100001000",
                      66 when "00110100001001",
                      66 when "00110100001010",
                      66 when "00110100001011",
                      66 when "00110100001100",
                      66 when "00110100001101",
                      66 when "00110100001110",
                      66 when "00110100001111",
                      66 when "00110100010000",
                      66 when "00110100010001",
                      66 when "00110100010010",
                      66 when "00110100010011",
                      66 when "00110100010100",
                      66 when "00110100010101",
                      66 when "00110100010110",
                      66 when "00110100010111",
                      66 when "00110100011000",
                      66 when "00110100011001",
                      66 when "00110100011010",
                      65 when "00110100011011",
                      65 when "00110100011100",
                      65 when "00110100011101",
                      65 when "00110100011110",
                      65 when "00110100011111",
                      65 when "00110100100000",
                      65 when "00110100100001",
                      65 when "00110100100010",
                      65 when "00110100100011",
                      65 when "00110100100100",
                      65 when "00110100100101",
                      65 when "00110100100110",
                      65 when "00110100100111",
                      65 when "00110100101000",
                      65 when "00110100101001",
                      65 when "00110100101010",
                      65 when "00110100101011",
                      65 when "00110100101100",
                      65 when "00110100101101",
                      65 when "00110100101110",
                      65 when "00110100101111",
                      65 when "00110100110000",
                      65 when "00110100110001",
                      65 when "00110100110010",
                      65 when "00110100110011",
                      65 when "00110100110100",
                      65 when "00110100110101",
                      65 when "00110100110110",
                      65 when "00110100110111",
                      65 when "00110100111000",
                      65 when "00110100111001",
                      65 when "00110100111010",
                      65 when "00110100111011",
                      65 when "00110100111100",
                      65 when "00110100111101",
                      65 when "00110100111110",
                      65 when "00110100111111",
                      65 when "00110101000000",
                      65 when "00110101000001",
                      65 when "00110101000010",
                      65 when "00110101000011",
                      65 when "00110101000100",
                      65 when "00110101000101",
                      65 when "00110101000110",
                      65 when "00110101000111",
                      65 when "00110101001000",
                      65 when "00110101001001",
                      65 when "00110101001010",
                      65 when "00110101001011",
                      65 when "00110101001100",
                      65 when "00110101001101",
                      65 when "00110101001110",
                      64 when "00110101001111",
                      64 when "00110101010000",
                      64 when "00110101010001",
                      64 when "00110101010010",
                      64 when "00110101010011",
                      64 when "00110101010100",
                      64 when "00110101010101",
                      64 when "00110101010110",
                      64 when "00110101010111",
                      64 when "00110101011000",
                      64 when "00110101011001",
                      64 when "00110101011010",
                      64 when "00110101011011",
                      64 when "00110101011100",
                      64 when "00110101011101",
                      64 when "00110101011110",
                      64 when "00110101011111",
                      64 when "00110101100000",
                      64 when "00110101100001",
                      64 when "00110101100010",
                      64 when "00110101100011",
                      64 when "00110101100100",
                      64 when "00110101100101",
                      64 when "00110101100110",
                      64 when "00110101100111",
                      64 when "00110101101000",
                      64 when "00110101101001",
                      64 when "00110101101010",
                      64 when "00110101101011",
                      64 when "00110101101100",
                      64 when "00110101101101",
                      64 when "00110101101110",
                      64 when "00110101101111",
                      64 when "00110101110000",
                      64 when "00110101110001",
                      64 when "00110101110010",
                      64 when "00110101110011",
                      64 when "00110101110100",
                      64 when "00110101110101",
                      64 when "00110101110110",
                      64 when "00110101110111",
                      64 when "00110101111000",
                      64 when "00110101111001",
                      64 when "00110101111010",
                      64 when "00110101111011",
                      64 when "00110101111100",
                      64 when "00110101111101",
                      64 when "00110101111110",
                      64 when "00110101111111",
                      64 when "00110110000000",
                      64 when "00110110000001",
                      64 when "00110110000010",
                      64 when "00110110000011",
                      64 when "00110110000100",
                      63 when "00110110000101",
                      63 when "00110110000110",
                      63 when "00110110000111",
                      63 when "00110110001000",
                      63 when "00110110001001",
                      63 when "00110110001010",
                      63 when "00110110001011",
                      63 when "00110110001100",
                      63 when "00110110001101",
                      63 when "00110110001110",
                      63 when "00110110001111",
                      63 when "00110110010000",
                      63 when "00110110010001",
                      63 when "00110110010010",
                      63 when "00110110010011",
                      63 when "00110110010100",
                      63 when "00110110010101",
                      63 when "00110110010110",
                      63 when "00110110010111",
                      63 when "00110110011000",
                      63 when "00110110011001",
                      63 when "00110110011010",
                      63 when "00110110011011",
                      63 when "00110110011100",
                      63 when "00110110011101",
                      63 when "00110110011110",
                      63 when "00110110011111",
                      63 when "00110110100000",
                      63 when "00110110100001",
                      63 when "00110110100010",
                      63 when "00110110100011",
                      63 when "00110110100100",
                      63 when "00110110100101",
                      63 when "00110110100110",
                      63 when "00110110100111",
                      63 when "00110110101000",
                      63 when "00110110101001",
                      63 when "00110110101010",
                      63 when "00110110101011",
                      63 when "00110110101100",
                      63 when "00110110101101",
                      63 when "00110110101110",
                      63 when "00110110101111",
                      63 when "00110110110000",
                      63 when "00110110110001",
                      63 when "00110110110010",
                      63 when "00110110110011",
                      63 when "00110110110100",
                      63 when "00110110110101",
                      63 when "00110110110110",
                      63 when "00110110110111",
                      63 when "00110110111000",
                      63 when "00110110111001",
                      63 when "00110110111010",
                      63 when "00110110111011",
                      62 when "00110110111100",
                      62 when "00110110111101",
                      62 when "00110110111110",
                      62 when "00110110111111",
                      62 when "00110111000000",
                      62 when "00110111000001",
                      62 when "00110111000010",
                      62 when "00110111000011",
                      62 when "00110111000100",
                      62 when "00110111000101",
                      62 when "00110111000110",
                      62 when "00110111000111",
                      62 when "00110111001000",
                      62 when "00110111001001",
                      62 when "00110111001010",
                      62 when "00110111001011",
                      62 when "00110111001100",
                      62 when "00110111001101",
                      62 when "00110111001110",
                      62 when "00110111001111",
                      62 when "00110111010000",
                      62 when "00110111010001",
                      62 when "00110111010010",
                      62 when "00110111010011",
                      62 when "00110111010100",
                      62 when "00110111010101",
                      62 when "00110111010110",
                      62 when "00110111010111",
                      62 when "00110111011000",
                      62 when "00110111011001",
                      62 when "00110111011010",
                      62 when "00110111011011",
                      62 when "00110111011100",
                      62 when "00110111011101",
                      62 when "00110111011110",
                      62 when "00110111011111",
                      62 when "00110111100000",
                      62 when "00110111100001",
                      62 when "00110111100010",
                      62 when "00110111100011",
                      62 when "00110111100100",
                      62 when "00110111100101",
                      62 when "00110111100110",
                      62 when "00110111100111",
                      62 when "00110111101000",
                      62 when "00110111101001",
                      62 when "00110111101010",
                      62 when "00110111101011",
                      62 when "00110111101100",
                      62 when "00110111101101",
                      62 when "00110111101110",
                      62 when "00110111101111",
                      62 when "00110111110000",
                      62 when "00110111110001",
                      62 when "00110111110010",
                      62 when "00110111110011",
                      62 when "00110111110100",
                      61 when "00110111110101",
                      61 when "00110111110110",
                      61 when "00110111110111",
                      61 when "00110111111000",
                      61 when "00110111111001",
                      61 when "00110111111010",
                      61 when "00110111111011",
                      61 when "00110111111100",
                      61 when "00110111111101",
                      61 when "00110111111110",
                      61 when "00110111111111",
                      61 when "00111000000000",
                      61 when "00111000000001",
                      61 when "00111000000010",
                      61 when "00111000000011",
                      61 when "00111000000100",
                      61 when "00111000000101",
                      61 when "00111000000110",
                      61 when "00111000000111",
                      61 when "00111000001000",
                      61 when "00111000001001",
                      61 when "00111000001010",
                      61 when "00111000001011",
                      61 when "00111000001100",
                      61 when "00111000001101",
                      61 when "00111000001110",
                      61 when "00111000001111",
                      61 when "00111000010000",
                      61 when "00111000010001",
                      61 when "00111000010010",
                      61 when "00111000010011",
                      61 when "00111000010100",
                      61 when "00111000010101",
                      61 when "00111000010110",
                      61 when "00111000010111",
                      61 when "00111000011000",
                      61 when "00111000011001",
                      61 when "00111000011010",
                      61 when "00111000011011",
                      61 when "00111000011100",
                      61 when "00111000011101",
                      61 when "00111000011110",
                      61 when "00111000011111",
                      61 when "00111000100000",
                      61 when "00111000100001",
                      61 when "00111000100010",
                      61 when "00111000100011",
                      61 when "00111000100100",
                      61 when "00111000100101",
                      61 when "00111000100110",
                      61 when "00111000100111",
                      61 when "00111000101000",
                      61 when "00111000101001",
                      61 when "00111000101010",
                      61 when "00111000101011",
                      61 when "00111000101100",
                      61 when "00111000101101",
                      61 when "00111000101110",
                      61 when "00111000101111",
                      60 when "00111000110000",
                      60 when "00111000110001",
                      60 when "00111000110010",
                      60 when "00111000110011",
                      60 when "00111000110100",
                      60 when "00111000110101",
                      60 when "00111000110110",
                      60 when "00111000110111",
                      60 when "00111000111000",
                      60 when "00111000111001",
                      60 when "00111000111010",
                      60 when "00111000111011",
                      60 when "00111000111100",
                      60 when "00111000111101",
                      60 when "00111000111110",
                      60 when "00111000111111",
                      60 when "00111001000000",
                      60 when "00111001000001",
                      60 when "00111001000010",
                      60 when "00111001000011",
                      60 when "00111001000100",
                      60 when "00111001000101",
                      60 when "00111001000110",
                      60 when "00111001000111",
                      60 when "00111001001000",
                      60 when "00111001001001",
                      60 when "00111001001010",
                      60 when "00111001001011",
                      60 when "00111001001100",
                      60 when "00111001001101",
                      60 when "00111001001110",
                      60 when "00111001001111",
                      60 when "00111001010000",
                      60 when "00111001010001",
                      60 when "00111001010010",
                      60 when "00111001010011",
                      60 when "00111001010100",
                      60 when "00111001010101",
                      60 when "00111001010110",
                      60 when "00111001010111",
                      60 when "00111001011000",
                      60 when "00111001011001",
                      60 when "00111001011010",
                      60 when "00111001011011",
                      60 when "00111001011100",
                      60 when "00111001011101",
                      60 when "00111001011110",
                      60 when "00111001011111",
                      60 when "00111001100000",
                      60 when "00111001100001",
                      60 when "00111001100010",
                      60 when "00111001100011",
                      60 when "00111001100100",
                      60 when "00111001100101",
                      60 when "00111001100110",
                      60 when "00111001100111",
                      60 when "00111001101000",
                      60 when "00111001101001",
                      60 when "00111001101010",
                      60 when "00111001101011",
                      60 when "00111001101100",
                      59 when "00111001101101",
                      59 when "00111001101110",
                      59 when "00111001101111",
                      59 when "00111001110000",
                      59 when "00111001110001",
                      59 when "00111001110010",
                      59 when "00111001110011",
                      59 when "00111001110100",
                      59 when "00111001110101",
                      59 when "00111001110110",
                      59 when "00111001110111",
                      59 when "00111001111000",
                      59 when "00111001111001",
                      59 when "00111001111010",
                      59 when "00111001111011",
                      59 when "00111001111100",
                      59 when "00111001111101",
                      59 when "00111001111110",
                      59 when "00111001111111",
                      59 when "00111010000000",
                      59 when "00111010000001",
                      59 when "00111010000010",
                      59 when "00111010000011",
                      59 when "00111010000100",
                      59 when "00111010000101",
                      59 when "00111010000110",
                      59 when "00111010000111",
                      59 when "00111010001000",
                      59 when "00111010001001",
                      59 when "00111010001010",
                      59 when "00111010001011",
                      59 when "00111010001100",
                      59 when "00111010001101",
                      59 when "00111010001110",
                      59 when "00111010001111",
                      59 when "00111010010000",
                      59 when "00111010010001",
                      59 when "00111010010010",
                      59 when "00111010010011",
                      59 when "00111010010100",
                      59 when "00111010010101",
                      59 when "00111010010110",
                      59 when "00111010010111",
                      59 when "00111010011000",
                      59 when "00111010011001",
                      59 when "00111010011010",
                      59 when "00111010011011",
                      59 when "00111010011100",
                      59 when "00111010011101",
                      59 when "00111010011110",
                      59 when "00111010011111",
                      59 when "00111010100000",
                      59 when "00111010100001",
                      59 when "00111010100010",
                      59 when "00111010100011",
                      59 when "00111010100100",
                      59 when "00111010100101",
                      59 when "00111010100110",
                      59 when "00111010100111",
                      59 when "00111010101000",
                      59 when "00111010101001",
                      59 when "00111010101010",
                      59 when "00111010101011",
                      59 when "00111010101100",
                      58 when "00111010101101",
                      58 when "00111010101110",
                      58 when "00111010101111",
                      58 when "00111010110000",
                      58 when "00111010110001",
                      58 when "00111010110010",
                      58 when "00111010110011",
                      58 when "00111010110100",
                      58 when "00111010110101",
                      58 when "00111010110110",
                      58 when "00111010110111",
                      58 when "00111010111000",
                      58 when "00111010111001",
                      58 when "00111010111010",
                      58 when "00111010111011",
                      58 when "00111010111100",
                      58 when "00111010111101",
                      58 when "00111010111110",
                      58 when "00111010111111",
                      58 when "00111011000000",
                      58 when "00111011000001",
                      58 when "00111011000010",
                      58 when "00111011000011",
                      58 when "00111011000100",
                      58 when "00111011000101",
                      58 when "00111011000110",
                      58 when "00111011000111",
                      58 when "00111011001000",
                      58 when "00111011001001",
                      58 when "00111011001010",
                      58 when "00111011001011",
                      58 when "00111011001100",
                      58 when "00111011001101",
                      58 when "00111011001110",
                      58 when "00111011001111",
                      58 when "00111011010000",
                      58 when "00111011010001",
                      58 when "00111011010010",
                      58 when "00111011010011",
                      58 when "00111011010100",
                      58 when "00111011010101",
                      58 when "00111011010110",
                      58 when "00111011010111",
                      58 when "00111011011000",
                      58 when "00111011011001",
                      58 when "00111011011010",
                      58 when "00111011011011",
                      58 when "00111011011100",
                      58 when "00111011011101",
                      58 when "00111011011110",
                      58 when "00111011011111",
                      58 when "00111011100000",
                      58 when "00111011100001",
                      58 when "00111011100010",
                      58 when "00111011100011",
                      58 when "00111011100100",
                      58 when "00111011100101",
                      58 when "00111011100110",
                      58 when "00111011100111",
                      58 when "00111011101000",
                      58 when "00111011101001",
                      58 when "00111011101010",
                      58 when "00111011101011",
                      58 when "00111011101100",
                      58 when "00111011101101",
                      57 when "00111011101110",
                      57 when "00111011101111",
                      57 when "00111011110000",
                      57 when "00111011110001",
                      57 when "00111011110010",
                      57 when "00111011110011",
                      57 when "00111011110100",
                      57 when "00111011110101",
                      57 when "00111011110110",
                      57 when "00111011110111",
                      57 when "00111011111000",
                      57 when "00111011111001",
                      57 when "00111011111010",
                      57 when "00111011111011",
                      57 when "00111011111100",
                      57 when "00111011111101",
                      57 when "00111011111110",
                      57 when "00111011111111",
                      57 when "00111100000000",
                      57 when "00111100000001",
                      57 when "00111100000010",
                      57 when "00111100000011",
                      57 when "00111100000100",
                      57 when "00111100000101",
                      57 when "00111100000110",
                      57 when "00111100000111",
                      57 when "00111100001000",
                      57 when "00111100001001",
                      57 when "00111100001010",
                      57 when "00111100001011",
                      57 when "00111100001100",
                      57 when "00111100001101",
                      57 when "00111100001110",
                      57 when "00111100001111",
                      57 when "00111100010000",
                      57 when "00111100010001",
                      57 when "00111100010010",
                      57 when "00111100010011",
                      57 when "00111100010100",
                      57 when "00111100010101",
                      57 when "00111100010110",
                      57 when "00111100010111",
                      57 when "00111100011000",
                      57 when "00111100011001",
                      57 when "00111100011010",
                      57 when "00111100011011",
                      57 when "00111100011100",
                      57 when "00111100011101",
                      57 when "00111100011110",
                      57 when "00111100011111",
                      57 when "00111100100000",
                      57 when "00111100100001",
                      57 when "00111100100010",
                      57 when "00111100100011",
                      57 when "00111100100100",
                      57 when "00111100100101",
                      57 when "00111100100110",
                      57 when "00111100100111",
                      57 when "00111100101000",
                      57 when "00111100101001",
                      57 when "00111100101010",
                      57 when "00111100101011",
                      57 when "00111100101100",
                      57 when "00111100101101",
                      57 when "00111100101110",
                      57 when "00111100101111",
                      57 when "00111100110000",
                      56 when "00111100110001",
                      56 when "00111100110010",
                      56 when "00111100110011",
                      56 when "00111100110100",
                      56 when "00111100110101",
                      56 when "00111100110110",
                      56 when "00111100110111",
                      56 when "00111100111000",
                      56 when "00111100111001",
                      56 when "00111100111010",
                      56 when "00111100111011",
                      56 when "00111100111100",
                      56 when "00111100111101",
                      56 when "00111100111110",
                      56 when "00111100111111",
                      56 when "00111101000000",
                      56 when "00111101000001",
                      56 when "00111101000010",
                      56 when "00111101000011",
                      56 when "00111101000100",
                      56 when "00111101000101",
                      56 when "00111101000110",
                      56 when "00111101000111",
                      56 when "00111101001000",
                      56 when "00111101001001",
                      56 when "00111101001010",
                      56 when "00111101001011",
                      56 when "00111101001100",
                      56 when "00111101001101",
                      56 when "00111101001110",
                      56 when "00111101001111",
                      56 when "00111101010000",
                      56 when "00111101010001",
                      56 when "00111101010010",
                      56 when "00111101010011",
                      56 when "00111101010100",
                      56 when "00111101010101",
                      56 when "00111101010110",
                      56 when "00111101010111",
                      56 when "00111101011000",
                      56 when "00111101011001",
                      56 when "00111101011010",
                      56 when "00111101011011",
                      56 when "00111101011100",
                      56 when "00111101011101",
                      56 when "00111101011110",
                      56 when "00111101011111",
                      56 when "00111101100000",
                      56 when "00111101100001",
                      56 when "00111101100010",
                      56 when "00111101100011",
                      56 when "00111101100100",
                      56 when "00111101100101",
                      56 when "00111101100110",
                      56 when "00111101100111",
                      56 when "00111101101000",
                      56 when "00111101101001",
                      56 when "00111101101010",
                      56 when "00111101101011",
                      56 when "00111101101100",
                      56 when "00111101101101",
                      56 when "00111101101110",
                      56 when "00111101101111",
                      56 when "00111101110000",
                      56 when "00111101110001",
                      56 when "00111101110010",
                      56 when "00111101110011",
                      56 when "00111101110100",
                      56 when "00111101110101",
                      56 when "00111101110110",
                      56 when "00111101110111",
                      55 when "00111101111000",
                      55 when "00111101111001",
                      55 when "00111101111010",
                      55 when "00111101111011",
                      55 when "00111101111100",
                      55 when "00111101111101",
                      55 when "00111101111110",
                      55 when "00111101111111",
                      55 when "00111110000000",
                      55 when "00111110000001",
                      55 when "00111110000010",
                      55 when "00111110000011",
                      55 when "00111110000100",
                      55 when "00111110000101",
                      55 when "00111110000110",
                      55 when "00111110000111",
                      55 when "00111110001000",
                      55 when "00111110001001",
                      55 when "00111110001010",
                      55 when "00111110001011",
                      55 when "00111110001100",
                      55 when "00111110001101",
                      55 when "00111110001110",
                      55 when "00111110001111",
                      55 when "00111110010000",
                      55 when "00111110010001",
                      55 when "00111110010010",
                      55 when "00111110010011",
                      55 when "00111110010100",
                      55 when "00111110010101",
                      55 when "00111110010110",
                      55 when "00111110010111",
                      55 when "00111110011000",
                      55 when "00111110011001",
                      55 when "00111110011010",
                      55 when "00111110011011",
                      55 when "00111110011100",
                      55 when "00111110011101",
                      55 when "00111110011110",
                      55 when "00111110011111",
                      55 when "00111110100000",
                      55 when "00111110100001",
                      55 when "00111110100010",
                      55 when "00111110100011",
                      55 when "00111110100100",
                      55 when "00111110100101",
                      55 when "00111110100110",
                      55 when "00111110100111",
                      55 when "00111110101000",
                      55 when "00111110101001",
                      55 when "00111110101010",
                      55 when "00111110101011",
                      55 when "00111110101100",
                      55 when "00111110101101",
                      55 when "00111110101110",
                      55 when "00111110101111",
                      55 when "00111110110000",
                      55 when "00111110110001",
                      55 when "00111110110010",
                      55 when "00111110110011",
                      55 when "00111110110100",
                      55 when "00111110110101",
                      55 when "00111110110110",
                      55 when "00111110110111",
                      55 when "00111110111000",
                      55 when "00111110111001",
                      55 when "00111110111010",
                      55 when "00111110111011",
                      55 when "00111110111100",
                      55 when "00111110111101",
                      55 when "00111110111110",
                      55 when "00111110111111",
                      54 when "00111111000000",
                      54 when "00111111000001",
                      54 when "00111111000010",
                      54 when "00111111000011",
                      54 when "00111111000100",
                      54 when "00111111000101",
                      54 when "00111111000110",
                      54 when "00111111000111",
                      54 when "00111111001000",
                      54 when "00111111001001",
                      54 when "00111111001010",
                      54 when "00111111001011",
                      54 when "00111111001100",
                      54 when "00111111001101",
                      54 when "00111111001110",
                      54 when "00111111001111",
                      54 when "00111111010000",
                      54 when "00111111010001",
                      54 when "00111111010010",
                      54 when "00111111010011",
                      54 when "00111111010100",
                      54 when "00111111010101",
                      54 when "00111111010110",
                      54 when "00111111010111",
                      54 when "00111111011000",
                      54 when "00111111011001",
                      54 when "00111111011010",
                      54 when "00111111011011",
                      54 when "00111111011100",
                      54 when "00111111011101",
                      54 when "00111111011110",
                      54 when "00111111011111",
                      54 when "00111111100000",
                      54 when "00111111100001",
                      54 when "00111111100010",
                      54 when "00111111100011",
                      54 when "00111111100100",
                      54 when "00111111100101",
                      54 when "00111111100110",
                      54 when "00111111100111",
                      54 when "00111111101000",
                      54 when "00111111101001",
                      54 when "00111111101010",
                      54 when "00111111101011",
                      54 when "00111111101100",
                      54 when "00111111101101",
                      54 when "00111111101110",
                      54 when "00111111101111",
                      54 when "00111111110000",
                      54 when "00111111110001",
                      54 when "00111111110010",
                      54 when "00111111110011",
                      54 when "00111111110100",
                      54 when "00111111110101",
                      54 when "00111111110110",
                      54 when "00111111110111",
                      54 when "00111111111000",
                      54 when "00111111111001",
                      54 when "00111111111010",
                      54 when "00111111111011",
                      54 when "00111111111100",
                      54 when "00111111111101",
                      54 when "00111111111110",
                      54 when "00111111111111",
                      54 when "01000000000000",
                      54 when "01000000000001",
                      54 when "01000000000010",
                      54 when "01000000000011",
                      54 when "01000000000100",
                      54 when "01000000000101",
                      54 when "01000000000110",
                      54 when "01000000000111",
                      54 when "01000000001000",
                      54 when "01000000001001",
                      54 when "01000000001010",
                      54 when "01000000001011",
                      53 when "01000000001100",
                      53 when "01000000001101",
                      53 when "01000000001110",
                      53 when "01000000001111",
                      53 when "01000000010000",
                      53 when "01000000010001",
                      53 when "01000000010010",
                      53 when "01000000010011",
                      53 when "01000000010100",
                      53 when "01000000010101",
                      53 when "01000000010110",
                      53 when "01000000010111",
                      53 when "01000000011000",
                      53 when "01000000011001",
                      53 when "01000000011010",
                      53 when "01000000011011",
                      53 when "01000000011100",
                      53 when "01000000011101",
                      53 when "01000000011110",
                      53 when "01000000011111",
                      53 when "01000000100000",
                      53 when "01000000100001",
                      53 when "01000000100010",
                      53 when "01000000100011",
                      53 when "01000000100100",
                      53 when "01000000100101",
                      53 when "01000000100110",
                      53 when "01000000100111",
                      53 when "01000000101000",
                      53 when "01000000101001",
                      53 when "01000000101010",
                      53 when "01000000101011",
                      53 when "01000000101100",
                      53 when "01000000101101",
                      53 when "01000000101110",
                      53 when "01000000101111",
                      53 when "01000000110000",
                      53 when "01000000110001",
                      53 when "01000000110010",
                      53 when "01000000110011",
                      53 when "01000000110100",
                      53 when "01000000110101",
                      53 when "01000000110110",
                      53 when "01000000110111",
                      53 when "01000000111000",
                      53 when "01000000111001",
                      53 when "01000000111010",
                      53 when "01000000111011",
                      53 when "01000000111100",
                      53 when "01000000111101",
                      53 when "01000000111110",
                      53 when "01000000111111",
                      53 when "01000001000000",
                      53 when "01000001000001",
                      53 when "01000001000010",
                      53 when "01000001000011",
                      53 when "01000001000100",
                      53 when "01000001000101",
                      53 when "01000001000110",
                      53 when "01000001000111",
                      53 when "01000001001000",
                      53 when "01000001001001",
                      53 when "01000001001010",
                      53 when "01000001001011",
                      53 when "01000001001100",
                      53 when "01000001001101",
                      53 when "01000001001110",
                      53 when "01000001001111",
                      53 when "01000001010000",
                      53 when "01000001010001",
                      53 when "01000001010010",
                      53 when "01000001010011",
                      53 when "01000001010100",
                      53 when "01000001010101",
                      53 when "01000001010110",
                      53 when "01000001010111",
                      53 when "01000001011000",
                      53 when "01000001011001",
                      52 when "01000001011010",
                      52 when "01000001011011",
                      52 when "01000001011100",
                      52 when "01000001011101",
                      52 when "01000001011110",
                      52 when "01000001011111",
                      52 when "01000001100000",
                      52 when "01000001100001",
                      52 when "01000001100010",
                      52 when "01000001100011",
                      52 when "01000001100100",
                      52 when "01000001100101",
                      52 when "01000001100110",
                      52 when "01000001100111",
                      52 when "01000001101000",
                      52 when "01000001101001",
                      52 when "01000001101010",
                      52 when "01000001101011",
                      52 when "01000001101100",
                      52 when "01000001101101",
                      52 when "01000001101110",
                      52 when "01000001101111",
                      52 when "01000001110000",
                      52 when "01000001110001",
                      52 when "01000001110010",
                      52 when "01000001110011",
                      52 when "01000001110100",
                      52 when "01000001110101",
                      52 when "01000001110110",
                      52 when "01000001110111",
                      52 when "01000001111000",
                      52 when "01000001111001",
                      52 when "01000001111010",
                      52 when "01000001111011",
                      52 when "01000001111100",
                      52 when "01000001111101",
                      52 when "01000001111110",
                      52 when "01000001111111",
                      52 when "01000010000000",
                      52 when "01000010000001",
                      52 when "01000010000010",
                      52 when "01000010000011",
                      52 when "01000010000100",
                      52 when "01000010000101",
                      52 when "01000010000110",
                      52 when "01000010000111",
                      52 when "01000010001000",
                      52 when "01000010001001",
                      52 when "01000010001010",
                      52 when "01000010001011",
                      52 when "01000010001100",
                      52 when "01000010001101",
                      52 when "01000010001110",
                      52 when "01000010001111",
                      52 when "01000010010000",
                      52 when "01000010010001",
                      52 when "01000010010010",
                      52 when "01000010010011",
                      52 when "01000010010100",
                      52 when "01000010010101",
                      52 when "01000010010110",
                      52 when "01000010010111",
                      52 when "01000010011000",
                      52 when "01000010011001",
                      52 when "01000010011010",
                      52 when "01000010011011",
                      52 when "01000010011100",
                      52 when "01000010011101",
                      52 when "01000010011110",
                      52 when "01000010011111",
                      52 when "01000010100000",
                      52 when "01000010100001",
                      52 when "01000010100010",
                      52 when "01000010100011",
                      52 when "01000010100100",
                      52 when "01000010100101",
                      52 when "01000010100110",
                      52 when "01000010100111",
                      52 when "01000010101000",
                      52 when "01000010101001",
                      52 when "01000010101010",
                      51 when "01000010101011",
                      51 when "01000010101100",
                      51 when "01000010101101",
                      51 when "01000010101110",
                      51 when "01000010101111",
                      51 when "01000010110000",
                      51 when "01000010110001",
                      51 when "01000010110010",
                      51 when "01000010110011",
                      51 when "01000010110100",
                      51 when "01000010110101",
                      51 when "01000010110110",
                      51 when "01000010110111",
                      51 when "01000010111000",
                      51 when "01000010111001",
                      51 when "01000010111010",
                      51 when "01000010111011",
                      51 when "01000010111100",
                      51 when "01000010111101",
                      51 when "01000010111110",
                      51 when "01000010111111",
                      51 when "01000011000000",
                      51 when "01000011000001",
                      51 when "01000011000010",
                      51 when "01000011000011",
                      51 when "01000011000100",
                      51 when "01000011000101",
                      51 when "01000011000110",
                      51 when "01000011000111",
                      51 when "01000011001000",
                      51 when "01000011001001",
                      51 when "01000011001010",
                      51 when "01000011001011",
                      51 when "01000011001100",
                      51 when "01000011001101",
                      51 when "01000011001110",
                      51 when "01000011001111",
                      51 when "01000011010000",
                      51 when "01000011010001",
                      51 when "01000011010010",
                      51 when "01000011010011",
                      51 when "01000011010100",
                      51 when "01000011010101",
                      51 when "01000011010110",
                      51 when "01000011010111",
                      51 when "01000011011000",
                      51 when "01000011011001",
                      51 when "01000011011010",
                      51 when "01000011011011",
                      51 when "01000011011100",
                      51 when "01000011011101",
                      51 when "01000011011110",
                      51 when "01000011011111",
                      51 when "01000011100000",
                      51 when "01000011100001",
                      51 when "01000011100010",
                      51 when "01000011100011",
                      51 when "01000011100100",
                      51 when "01000011100101",
                      51 when "01000011100110",
                      51 when "01000011100111",
                      51 when "01000011101000",
                      51 when "01000011101001",
                      51 when "01000011101010",
                      51 when "01000011101011",
                      51 when "01000011101100",
                      51 when "01000011101101",
                      51 when "01000011101110",
                      51 when "01000011101111",
                      51 when "01000011110000",
                      51 when "01000011110001",
                      51 when "01000011110010",
                      51 when "01000011110011",
                      51 when "01000011110100",
                      51 when "01000011110101",
                      51 when "01000011110110",
                      51 when "01000011110111",
                      51 when "01000011111000",
                      51 when "01000011111001",
                      51 when "01000011111010",
                      51 when "01000011111011",
                      51 when "01000011111100",
                      51 when "01000011111101",
                      51 when "01000011111110",
                      51 when "01000011111111",
                      50 when "01000100000000",
                      50 when "01000100000001",
                      50 when "01000100000010",
                      50 when "01000100000011",
                      50 when "01000100000100",
                      50 when "01000100000101",
                      50 when "01000100000110",
                      50 when "01000100000111",
                      50 when "01000100001000",
                      50 when "01000100001001",
                      50 when "01000100001010",
                      50 when "01000100001011",
                      50 when "01000100001100",
                      50 when "01000100001101",
                      50 when "01000100001110",
                      50 when "01000100001111",
                      50 when "01000100010000",
                      50 when "01000100010001",
                      50 when "01000100010010",
                      50 when "01000100010011",
                      50 when "01000100010100",
                      50 when "01000100010101",
                      50 when "01000100010110",
                      50 when "01000100010111",
                      50 when "01000100011000",
                      50 when "01000100011001",
                      50 when "01000100011010",
                      50 when "01000100011011",
                      50 when "01000100011100",
                      50 when "01000100011101",
                      50 when "01000100011110",
                      50 when "01000100011111",
                      50 when "01000100100000",
                      50 when "01000100100001",
                      50 when "01000100100010",
                      50 when "01000100100011",
                      50 when "01000100100100",
                      50 when "01000100100101",
                      50 when "01000100100110",
                      50 when "01000100100111",
                      50 when "01000100101000",
                      50 when "01000100101001",
                      50 when "01000100101010",
                      50 when "01000100101011",
                      50 when "01000100101100",
                      50 when "01000100101101",
                      50 when "01000100101110",
                      50 when "01000100101111",
                      50 when "01000100110000",
                      50 when "01000100110001",
                      50 when "01000100110010",
                      50 when "01000100110011",
                      50 when "01000100110100",
                      50 when "01000100110101",
                      50 when "01000100110110",
                      50 when "01000100110111",
                      50 when "01000100111000",
                      50 when "01000100111001",
                      50 when "01000100111010",
                      50 when "01000100111011",
                      50 when "01000100111100",
                      50 when "01000100111101",
                      50 when "01000100111110",
                      50 when "01000100111111",
                      50 when "01000101000000",
                      50 when "01000101000001",
                      50 when "01000101000010",
                      50 when "01000101000011",
                      50 when "01000101000100",
                      50 when "01000101000101",
                      50 when "01000101000110",
                      50 when "01000101000111",
                      50 when "01000101001000",
                      50 when "01000101001001",
                      50 when "01000101001010",
                      50 when "01000101001011",
                      50 when "01000101001100",
                      50 when "01000101001101",
                      50 when "01000101001110",
                      50 when "01000101001111",
                      50 when "01000101010000",
                      50 when "01000101010001",
                      50 when "01000101010010",
                      50 when "01000101010011",
                      50 when "01000101010100",
                      50 when "01000101010101",
                      50 when "01000101010110",
                      49 when "01000101010111",
                      49 when "01000101011000",
                      49 when "01000101011001",
                      49 when "01000101011010",
                      49 when "01000101011011",
                      49 when "01000101011100",
                      49 when "01000101011101",
                      49 when "01000101011110",
                      49 when "01000101011111",
                      49 when "01000101100000",
                      49 when "01000101100001",
                      49 when "01000101100010",
                      49 when "01000101100011",
                      49 when "01000101100100",
                      49 when "01000101100101",
                      49 when "01000101100110",
                      49 when "01000101100111",
                      49 when "01000101101000",
                      49 when "01000101101001",
                      49 when "01000101101010",
                      49 when "01000101101011",
                      49 when "01000101101100",
                      49 when "01000101101101",
                      49 when "01000101101110",
                      49 when "01000101101111",
                      49 when "01000101110000",
                      49 when "01000101110001",
                      49 when "01000101110010",
                      49 when "01000101110011",
                      49 when "01000101110100",
                      49 when "01000101110101",
                      49 when "01000101110110",
                      49 when "01000101110111",
                      49 when "01000101111000",
                      49 when "01000101111001",
                      49 when "01000101111010",
                      49 when "01000101111011",
                      49 when "01000101111100",
                      49 when "01000101111101",
                      49 when "01000101111110",
                      49 when "01000101111111",
                      49 when "01000110000000",
                      49 when "01000110000001",
                      49 when "01000110000010",
                      49 when "01000110000011",
                      49 when "01000110000100",
                      49 when "01000110000101",
                      49 when "01000110000110",
                      49 when "01000110000111",
                      49 when "01000110001000",
                      49 when "01000110001001",
                      49 when "01000110001010",
                      49 when "01000110001011",
                      49 when "01000110001100",
                      49 when "01000110001101",
                      49 when "01000110001110",
                      49 when "01000110001111",
                      49 when "01000110010000",
                      49 when "01000110010001",
                      49 when "01000110010010",
                      49 when "01000110010011",
                      49 when "01000110010100",
                      49 when "01000110010101",
                      49 when "01000110010110",
                      49 when "01000110010111",
                      49 when "01000110011000",
                      49 when "01000110011001",
                      49 when "01000110011010",
                      49 when "01000110011011",
                      49 when "01000110011100",
                      49 when "01000110011101",
                      49 when "01000110011110",
                      49 when "01000110011111",
                      49 when "01000110100000",
                      49 when "01000110100001",
                      49 when "01000110100010",
                      49 when "01000110100011",
                      49 when "01000110100100",
                      49 when "01000110100101",
                      49 when "01000110100110",
                      49 when "01000110100111",
                      49 when "01000110101000",
                      49 when "01000110101001",
                      49 when "01000110101010",
                      49 when "01000110101011",
                      49 when "01000110101100",
                      49 when "01000110101101",
                      49 when "01000110101110",
                      49 when "01000110101111",
                      49 when "01000110110000",
                      49 when "01000110110001",
                      49 when "01000110110010",
                      48 when "01000110110011",
                      48 when "01000110110100",
                      48 when "01000110110101",
                      48 when "01000110110110",
                      48 when "01000110110111",
                      48 when "01000110111000",
                      48 when "01000110111001",
                      48 when "01000110111010",
                      48 when "01000110111011",
                      48 when "01000110111100",
                      48 when "01000110111101",
                      48 when "01000110111110",
                      48 when "01000110111111",
                      48 when "01000111000000",
                      48 when "01000111000001",
                      48 when "01000111000010",
                      48 when "01000111000011",
                      48 when "01000111000100",
                      48 when "01000111000101",
                      48 when "01000111000110",
                      48 when "01000111000111",
                      48 when "01000111001000",
                      48 when "01000111001001",
                      48 when "01000111001010",
                      48 when "01000111001011",
                      48 when "01000111001100",
                      48 when "01000111001101",
                      48 when "01000111001110",
                      48 when "01000111001111",
                      48 when "01000111010000",
                      48 when "01000111010001",
                      48 when "01000111010010",
                      48 when "01000111010011",
                      48 when "01000111010100",
                      48 when "01000111010101",
                      48 when "01000111010110",
                      48 when "01000111010111",
                      48 when "01000111011000",
                      48 when "01000111011001",
                      48 when "01000111011010",
                      48 when "01000111011011",
                      48 when "01000111011100",
                      48 when "01000111011101",
                      48 when "01000111011110",
                      48 when "01000111011111",
                      48 when "01000111100000",
                      48 when "01000111100001",
                      48 when "01000111100010",
                      48 when "01000111100011",
                      48 when "01000111100100",
                      48 when "01000111100101",
                      48 when "01000111100110",
                      48 when "01000111100111",
                      48 when "01000111101000",
                      48 when "01000111101001",
                      48 when "01000111101010",
                      48 when "01000111101011",
                      48 when "01000111101100",
                      48 when "01000111101101",
                      48 when "01000111101110",
                      48 when "01000111101111",
                      48 when "01000111110000",
                      48 when "01000111110001",
                      48 when "01000111110010",
                      48 when "01000111110011",
                      48 when "01000111110100",
                      48 when "01000111110101",
                      48 when "01000111110110",
                      48 when "01000111110111",
                      48 when "01000111111000",
                      48 when "01000111111001",
                      48 when "01000111111010",
                      48 when "01000111111011",
                      48 when "01000111111100",
                      48 when "01000111111101",
                      48 when "01000111111110",
                      48 when "01000111111111",
                      48 when "01001000000000",
                      48 when "01001000000001",
                      48 when "01001000000010",
                      48 when "01001000000011",
                      48 when "01001000000100",
                      48 when "01001000000101",
                      48 when "01001000000110",
                      48 when "01001000000111",
                      48 when "01001000001000",
                      48 when "01001000001001",
                      48 when "01001000001010",
                      48 when "01001000001011",
                      48 when "01001000001100",
                      48 when "01001000001101",
                      48 when "01001000001110",
                      48 when "01001000001111",
                      48 when "01001000010000",
                      48 when "01001000010001",
                      47 when "01001000010010",
                      47 when "01001000010011",
                      47 when "01001000010100",
                      47 when "01001000010101",
                      47 when "01001000010110",
                      47 when "01001000010111",
                      47 when "01001000011000",
                      47 when "01001000011001",
                      47 when "01001000011010",
                      47 when "01001000011011",
                      47 when "01001000011100",
                      47 when "01001000011101",
                      47 when "01001000011110",
                      47 when "01001000011111",
                      47 when "01001000100000",
                      47 when "01001000100001",
                      47 when "01001000100010",
                      47 when "01001000100011",
                      47 when "01001000100100",
                      47 when "01001000100101",
                      47 when "01001000100110",
                      47 when "01001000100111",
                      47 when "01001000101000",
                      47 when "01001000101001",
                      47 when "01001000101010",
                      47 when "01001000101011",
                      47 when "01001000101100",
                      47 when "01001000101101",
                      47 when "01001000101110",
                      47 when "01001000101111",
                      47 when "01001000110000",
                      47 when "01001000110001",
                      47 when "01001000110010",
                      47 when "01001000110011",
                      47 when "01001000110100",
                      47 when "01001000110101",
                      47 when "01001000110110",
                      47 when "01001000110111",
                      47 when "01001000111000",
                      47 when "01001000111001",
                      47 when "01001000111010",
                      47 when "01001000111011",
                      47 when "01001000111100",
                      47 when "01001000111101",
                      47 when "01001000111110",
                      47 when "01001000111111",
                      47 when "01001001000000",
                      47 when "01001001000001",
                      47 when "01001001000010",
                      47 when "01001001000011",
                      47 when "01001001000100",
                      47 when "01001001000101",
                      47 when "01001001000110",
                      47 when "01001001000111",
                      47 when "01001001001000",
                      47 when "01001001001001",
                      47 when "01001001001010",
                      47 when "01001001001011",
                      47 when "01001001001100",
                      47 when "01001001001101",
                      47 when "01001001001110",
                      47 when "01001001001111",
                      47 when "01001001010000",
                      47 when "01001001010001",
                      47 when "01001001010010",
                      47 when "01001001010011",
                      47 when "01001001010100",
                      47 when "01001001010101",
                      47 when "01001001010110",
                      47 when "01001001010111",
                      47 when "01001001011000",
                      47 when "01001001011001",
                      47 when "01001001011010",
                      47 when "01001001011011",
                      47 when "01001001011100",
                      47 when "01001001011101",
                      47 when "01001001011110",
                      47 when "01001001011111",
                      47 when "01001001100000",
                      47 when "01001001100001",
                      47 when "01001001100010",
                      47 when "01001001100011",
                      47 when "01001001100100",
                      47 when "01001001100101",
                      47 when "01001001100110",
                      47 when "01001001100111",
                      47 when "01001001101000",
                      47 when "01001001101001",
                      47 when "01001001101010",
                      47 when "01001001101011",
                      47 when "01001001101100",
                      47 when "01001001101101",
                      47 when "01001001101110",
                      47 when "01001001101111",
                      47 when "01001001110000",
                      47 when "01001001110001",
                      47 when "01001001110010",
                      47 when "01001001110011",
                      47 when "01001001110100",
                      47 when "01001001110101",
                      46 when "01001001110110",
                      46 when "01001001110111",
                      46 when "01001001111000",
                      46 when "01001001111001",
                      46 when "01001001111010",
                      46 when "01001001111011",
                      46 when "01001001111100",
                      46 when "01001001111101",
                      46 when "01001001111110",
                      46 when "01001001111111",
                      46 when "01001010000000",
                      46 when "01001010000001",
                      46 when "01001010000010",
                      46 when "01001010000011",
                      46 when "01001010000100",
                      46 when "01001010000101",
                      46 when "01001010000110",
                      46 when "01001010000111",
                      46 when "01001010001000",
                      46 when "01001010001001",
                      46 when "01001010001010",
                      46 when "01001010001011",
                      46 when "01001010001100",
                      46 when "01001010001101",
                      46 when "01001010001110",
                      46 when "01001010001111",
                      46 when "01001010010000",
                      46 when "01001010010001",
                      46 when "01001010010010",
                      46 when "01001010010011",
                      46 when "01001010010100",
                      46 when "01001010010101",
                      46 when "01001010010110",
                      46 when "01001010010111",
                      46 when "01001010011000",
                      46 when "01001010011001",
                      46 when "01001010011010",
                      46 when "01001010011011",
                      46 when "01001010011100",
                      46 when "01001010011101",
                      46 when "01001010011110",
                      46 when "01001010011111",
                      46 when "01001010100000",
                      46 when "01001010100001",
                      46 when "01001010100010",
                      46 when "01001010100011",
                      46 when "01001010100100",
                      46 when "01001010100101",
                      46 when "01001010100110",
                      46 when "01001010100111",
                      46 when "01001010101000",
                      46 when "01001010101001",
                      46 when "01001010101010",
                      46 when "01001010101011",
                      46 when "01001010101100",
                      46 when "01001010101101",
                      46 when "01001010101110",
                      46 when "01001010101111",
                      46 when "01001010110000",
                      46 when "01001010110001",
                      46 when "01001010110010",
                      46 when "01001010110011",
                      46 when "01001010110100",
                      46 when "01001010110101",
                      46 when "01001010110110",
                      46 when "01001010110111",
                      46 when "01001010111000",
                      46 when "01001010111001",
                      46 when "01001010111010",
                      46 when "01001010111011",
                      46 when "01001010111100",
                      46 when "01001010111101",
                      46 when "01001010111110",
                      46 when "01001010111111",
                      46 when "01001011000000",
                      46 when "01001011000001",
                      46 when "01001011000010",
                      46 when "01001011000011",
                      46 when "01001011000100",
                      46 when "01001011000101",
                      46 when "01001011000110",
                      46 when "01001011000111",
                      46 when "01001011001000",
                      46 when "01001011001001",
                      46 when "01001011001010",
                      46 when "01001011001011",
                      46 when "01001011001100",
                      46 when "01001011001101",
                      46 when "01001011001110",
                      46 when "01001011001111",
                      46 when "01001011010000",
                      46 when "01001011010001",
                      46 when "01001011010010",
                      46 when "01001011010011",
                      46 when "01001011010100",
                      46 when "01001011010101",
                      46 when "01001011010110",
                      46 when "01001011010111",
                      46 when "01001011011000",
                      46 when "01001011011001",
                      46 when "01001011011010",
                      46 when "01001011011011",
                      46 when "01001011011100",
                      46 when "01001011011101",
                      45 when "01001011011110",
                      45 when "01001011011111",
                      45 when "01001011100000",
                      45 when "01001011100001",
                      45 when "01001011100010",
                      45 when "01001011100011",
                      45 when "01001011100100",
                      45 when "01001011100101",
                      45 when "01001011100110",
                      45 when "01001011100111",
                      45 when "01001011101000",
                      45 when "01001011101001",
                      45 when "01001011101010",
                      45 when "01001011101011",
                      45 when "01001011101100",
                      45 when "01001011101101",
                      45 when "01001011101110",
                      45 when "01001011101111",
                      45 when "01001011110000",
                      45 when "01001011110001",
                      45 when "01001011110010",
                      45 when "01001011110011",
                      45 when "01001011110100",
                      45 when "01001011110101",
                      45 when "01001011110110",
                      45 when "01001011110111",
                      45 when "01001011111000",
                      45 when "01001011111001",
                      45 when "01001011111010",
                      45 when "01001011111011",
                      45 when "01001011111100",
                      45 when "01001011111101",
                      45 when "01001011111110",
                      45 when "01001011111111",
                      45 when "01001100000000",
                      45 when "01001100000001",
                      45 when "01001100000010",
                      45 when "01001100000011",
                      45 when "01001100000100",
                      45 when "01001100000101",
                      45 when "01001100000110",
                      45 when "01001100000111",
                      45 when "01001100001000",
                      45 when "01001100001001",
                      45 when "01001100001010",
                      45 when "01001100001011",
                      45 when "01001100001100",
                      45 when "01001100001101",
                      45 when "01001100001110",
                      45 when "01001100001111",
                      45 when "01001100010000",
                      45 when "01001100010001",
                      45 when "01001100010010",
                      45 when "01001100010011",
                      45 when "01001100010100",
                      45 when "01001100010101",
                      45 when "01001100010110",
                      45 when "01001100010111",
                      45 when "01001100011000",
                      45 when "01001100011001",
                      45 when "01001100011010",
                      45 when "01001100011011",
                      45 when "01001100011100",
                      45 when "01001100011101",
                      45 when "01001100011110",
                      45 when "01001100011111",
                      45 when "01001100100000",
                      45 when "01001100100001",
                      45 when "01001100100010",
                      45 when "01001100100011",
                      45 when "01001100100100",
                      45 when "01001100100101",
                      45 when "01001100100110",
                      45 when "01001100100111",
                      45 when "01001100101000",
                      45 when "01001100101001",
                      45 when "01001100101010",
                      45 when "01001100101011",
                      45 when "01001100101100",
                      45 when "01001100101101",
                      45 when "01001100101110",
                      45 when "01001100101111",
                      45 when "01001100110000",
                      45 when "01001100110001",
                      45 when "01001100110010",
                      45 when "01001100110011",
                      45 when "01001100110100",
                      45 when "01001100110101",
                      45 when "01001100110110",
                      45 when "01001100110111",
                      45 when "01001100111000",
                      45 when "01001100111001",
                      45 when "01001100111010",
                      45 when "01001100111011",
                      45 when "01001100111100",
                      45 when "01001100111101",
                      45 when "01001100111110",
                      45 when "01001100111111",
                      45 when "01001101000000",
                      45 when "01001101000001",
                      45 when "01001101000010",
                      45 when "01001101000011",
                      45 when "01001101000100",
                      45 when "01001101000101",
                      45 when "01001101000110",
                      45 when "01001101000111",
                      45 when "01001101001000",
                      45 when "01001101001001",
                      44 when "01001101001010",
                      44 when "01001101001011",
                      44 when "01001101001100",
                      44 when "01001101001101",
                      44 when "01001101001110",
                      44 when "01001101001111",
                      44 when "01001101010000",
                      44 when "01001101010001",
                      44 when "01001101010010",
                      44 when "01001101010011",
                      44 when "01001101010100",
                      44 when "01001101010101",
                      44 when "01001101010110",
                      44 when "01001101010111",
                      44 when "01001101011000",
                      44 when "01001101011001",
                      44 when "01001101011010",
                      44 when "01001101011011",
                      44 when "01001101011100",
                      44 when "01001101011101",
                      44 when "01001101011110",
                      44 when "01001101011111",
                      44 when "01001101100000",
                      44 when "01001101100001",
                      44 when "01001101100010",
                      44 when "01001101100011",
                      44 when "01001101100100",
                      44 when "01001101100101",
                      44 when "01001101100110",
                      44 when "01001101100111",
                      44 when "01001101101000",
                      44 when "01001101101001",
                      44 when "01001101101010",
                      44 when "01001101101011",
                      44 when "01001101101100",
                      44 when "01001101101101",
                      44 when "01001101101110",
                      44 when "01001101101111",
                      44 when "01001101110000",
                      44 when "01001101110001",
                      44 when "01001101110010",
                      44 when "01001101110011",
                      44 when "01001101110100",
                      44 when "01001101110101",
                      44 when "01001101110110",
                      44 when "01001101110111",
                      44 when "01001101111000",
                      44 when "01001101111001",
                      44 when "01001101111010",
                      44 when "01001101111011",
                      44 when "01001101111100",
                      44 when "01001101111101",
                      44 when "01001101111110",
                      44 when "01001101111111",
                      44 when "01001110000000",
                      44 when "01001110000001",
                      44 when "01001110000010",
                      44 when "01001110000011",
                      44 when "01001110000100",
                      44 when "01001110000101",
                      44 when "01001110000110",
                      44 when "01001110000111",
                      44 when "01001110001000",
                      44 when "01001110001001",
                      44 when "01001110001010",
                      44 when "01001110001011",
                      44 when "01001110001100",
                      44 when "01001110001101",
                      44 when "01001110001110",
                      44 when "01001110001111",
                      44 when "01001110010000",
                      44 when "01001110010001",
                      44 when "01001110010010",
                      44 when "01001110010011",
                      44 when "01001110010100",
                      44 when "01001110010101",
                      44 when "01001110010110",
                      44 when "01001110010111",
                      44 when "01001110011000",
                      44 when "01001110011001",
                      44 when "01001110011010",
                      44 when "01001110011011",
                      44 when "01001110011100",
                      44 when "01001110011101",
                      44 when "01001110011110",
                      44 when "01001110011111",
                      44 when "01001110100000",
                      44 when "01001110100001",
                      44 when "01001110100010",
                      44 when "01001110100011",
                      44 when "01001110100100",
                      44 when "01001110100101",
                      44 when "01001110100110",
                      44 when "01001110100111",
                      44 when "01001110101000",
                      44 when "01001110101001",
                      44 when "01001110101010",
                      44 when "01001110101011",
                      44 when "01001110101100",
                      44 when "01001110101101",
                      44 when "01001110101110",
                      44 when "01001110101111",
                      44 when "01001110110000",
                      44 when "01001110110001",
                      44 when "01001110110010",
                      44 when "01001110110011",
                      44 when "01001110110100",
                      44 when "01001110110101",
                      44 when "01001110110110",
                      44 when "01001110110111",
                      44 when "01001110111000",
                      44 when "01001110111001",
                      44 when "01001110111010",
                      44 when "01001110111011",
                      43 when "01001110111100",
                      43 when "01001110111101",
                      43 when "01001110111110",
                      43 when "01001110111111",
                      43 when "01001111000000",
                      43 when "01001111000001",
                      43 when "01001111000010",
                      43 when "01001111000011",
                      43 when "01001111000100",
                      43 when "01001111000101",
                      43 when "01001111000110",
                      43 when "01001111000111",
                      43 when "01001111001000",
                      43 when "01001111001001",
                      43 when "01001111001010",
                      43 when "01001111001011",
                      43 when "01001111001100",
                      43 when "01001111001101",
                      43 when "01001111001110",
                      43 when "01001111001111",
                      43 when "01001111010000",
                      43 when "01001111010001",
                      43 when "01001111010010",
                      43 when "01001111010011",
                      43 when "01001111010100",
                      43 when "01001111010101",
                      43 when "01001111010110",
                      43 when "01001111010111",
                      43 when "01001111011000",
                      43 when "01001111011001",
                      43 when "01001111011010",
                      43 when "01001111011011",
                      43 when "01001111011100",
                      43 when "01001111011101",
                      43 when "01001111011110",
                      43 when "01001111011111",
                      43 when "01001111100000",
                      43 when "01001111100001",
                      43 when "01001111100010",
                      43 when "01001111100011",
                      43 when "01001111100100",
                      43 when "01001111100101",
                      43 when "01001111100110",
                      43 when "01001111100111",
                      43 when "01001111101000",
                      43 when "01001111101001",
                      43 when "01001111101010",
                      43 when "01001111101011",
                      43 when "01001111101100",
                      43 when "01001111101101",
                      43 when "01001111101110",
                      43 when "01001111101111",
                      43 when "01001111110000",
                      43 when "01001111110001",
                      43 when "01001111110010",
                      43 when "01001111110011",
                      43 when "01001111110100",
                      43 when "01001111110101",
                      43 when "01001111110110",
                      43 when "01001111110111",
                      43 when "01001111111000",
                      43 when "01001111111001",
                      43 when "01001111111010",
                      43 when "01001111111011",
                      43 when "01001111111100",
                      43 when "01001111111101",
                      43 when "01001111111110",
                      43 when "01001111111111",
                      43 when "01010000000000",
                      43 when "01010000000001",
                      43 when "01010000000010",
                      43 when "01010000000011",
                      43 when "01010000000100",
                      43 when "01010000000101",
                      43 when "01010000000110",
                      43 when "01010000000111",
                      43 when "01010000001000",
                      43 when "01010000001001",
                      43 when "01010000001010",
                      43 when "01010000001011",
                      43 when "01010000001100",
                      43 when "01010000001101",
                      43 when "01010000001110",
                      43 when "01010000001111",
                      43 when "01010000010000",
                      43 when "01010000010001",
                      43 when "01010000010010",
                      43 when "01010000010011",
                      43 when "01010000010100",
                      43 when "01010000010101",
                      43 when "01010000010110",
                      43 when "01010000010111",
                      43 when "01010000011000",
                      43 when "01010000011001",
                      43 when "01010000011010",
                      43 when "01010000011011",
                      43 when "01010000011100",
                      43 when "01010000011101",
                      43 when "01010000011110",
                      43 when "01010000011111",
                      43 when "01010000100000",
                      43 when "01010000100001",
                      43 when "01010000100010",
                      43 when "01010000100011",
                      43 when "01010000100100",
                      43 when "01010000100101",
                      43 when "01010000100110",
                      43 when "01010000100111",
                      43 when "01010000101000",
                      43 when "01010000101001",
                      43 when "01010000101010",
                      43 when "01010000101011",
                      43 when "01010000101100",
                      43 when "01010000101101",
                      43 when "01010000101110",
                      43 when "01010000101111",
                      43 when "01010000110000",
                      43 when "01010000110001",
                      43 when "01010000110010",
                      42 when "01010000110011",
                      42 when "01010000110100",
                      42 when "01010000110101",
                      42 when "01010000110110",
                      42 when "01010000110111",
                      42 when "01010000111000",
                      42 when "01010000111001",
                      42 when "01010000111010",
                      42 when "01010000111011",
                      42 when "01010000111100",
                      42 when "01010000111101",
                      42 when "01010000111110",
                      42 when "01010000111111",
                      42 when "01010001000000",
                      42 when "01010001000001",
                      42 when "01010001000010",
                      42 when "01010001000011",
                      42 when "01010001000100",
                      42 when "01010001000101",
                      42 when "01010001000110",
                      42 when "01010001000111",
                      42 when "01010001001000",
                      42 when "01010001001001",
                      42 when "01010001001010",
                      42 when "01010001001011",
                      42 when "01010001001100",
                      42 when "01010001001101",
                      42 when "01010001001110",
                      42 when "01010001001111",
                      42 when "01010001010000",
                      42 when "01010001010001",
                      42 when "01010001010010",
                      42 when "01010001010011",
                      42 when "01010001010100",
                      42 when "01010001010101",
                      42 when "01010001010110",
                      42 when "01010001010111",
                      42 when "01010001011000",
                      42 when "01010001011001",
                      42 when "01010001011010",
                      42 when "01010001011011",
                      42 when "01010001011100",
                      42 when "01010001011101",
                      42 when "01010001011110",
                      42 when "01010001011111",
                      42 when "01010001100000",
                      42 when "01010001100001",
                      42 when "01010001100010",
                      42 when "01010001100011",
                      42 when "01010001100100",
                      42 when "01010001100101",
                      42 when "01010001100110",
                      42 when "01010001100111",
                      42 when "01010001101000",
                      42 when "01010001101001",
                      42 when "01010001101010",
                      42 when "01010001101011",
                      42 when "01010001101100",
                      42 when "01010001101101",
                      42 when "01010001101110",
                      42 when "01010001101111",
                      42 when "01010001110000",
                      42 when "01010001110001",
                      42 when "01010001110010",
                      42 when "01010001110011",
                      42 when "01010001110100",
                      42 when "01010001110101",
                      42 when "01010001110110",
                      42 when "01010001110111",
                      42 when "01010001111000",
                      42 when "01010001111001",
                      42 when "01010001111010",
                      42 when "01010001111011",
                      42 when "01010001111100",
                      42 when "01010001111101",
                      42 when "01010001111110",
                      42 when "01010001111111",
                      42 when "01010010000000",
                      42 when "01010010000001",
                      42 when "01010010000010",
                      42 when "01010010000011",
                      42 when "01010010000100",
                      42 when "01010010000101",
                      42 when "01010010000110",
                      42 when "01010010000111",
                      42 when "01010010001000",
                      42 when "01010010001001",
                      42 when "01010010001010",
                      42 when "01010010001011",
                      42 when "01010010001100",
                      42 when "01010010001101",
                      42 when "01010010001110",
                      42 when "01010010001111",
                      42 when "01010010010000",
                      42 when "01010010010001",
                      42 when "01010010010010",
                      42 when "01010010010011",
                      42 when "01010010010100",
                      42 when "01010010010101",
                      42 when "01010010010110",
                      42 when "01010010010111",
                      42 when "01010010011000",
                      42 when "01010010011001",
                      42 when "01010010011010",
                      42 when "01010010011011",
                      42 when "01010010011100",
                      42 when "01010010011101",
                      42 when "01010010011110",
                      42 when "01010010011111",
                      42 when "01010010100000",
                      42 when "01010010100001",
                      42 when "01010010100010",
                      42 when "01010010100011",
                      42 when "01010010100100",
                      42 when "01010010100101",
                      42 when "01010010100110",
                      42 when "01010010100111",
                      42 when "01010010101000",
                      42 when "01010010101001",
                      42 when "01010010101010",
                      42 when "01010010101011",
                      42 when "01010010101100",
                      42 when "01010010101101",
                      42 when "01010010101110",
                      41 when "01010010101111",
                      41 when "01010010110000",
                      41 when "01010010110001",
                      41 when "01010010110010",
                      41 when "01010010110011",
                      41 when "01010010110100",
                      41 when "01010010110101",
                      41 when "01010010110110",
                      41 when "01010010110111",
                      41 when "01010010111000",
                      41 when "01010010111001",
                      41 when "01010010111010",
                      41 when "01010010111011",
                      41 when "01010010111100",
                      41 when "01010010111101",
                      41 when "01010010111110",
                      41 when "01010010111111",
                      41 when "01010011000000",
                      41 when "01010011000001",
                      41 when "01010011000010",
                      41 when "01010011000011",
                      41 when "01010011000100",
                      41 when "01010011000101",
                      41 when "01010011000110",
                      41 when "01010011000111",
                      41 when "01010011001000",
                      41 when "01010011001001",
                      41 when "01010011001010",
                      41 when "01010011001011",
                      41 when "01010011001100",
                      41 when "01010011001101",
                      41 when "01010011001110",
                      41 when "01010011001111",
                      41 when "01010011010000",
                      41 when "01010011010001",
                      41 when "01010011010010",
                      41 when "01010011010011",
                      41 when "01010011010100",
                      41 when "01010011010101",
                      41 when "01010011010110",
                      41 when "01010011010111",
                      41 when "01010011011000",
                      41 when "01010011011001",
                      41 when "01010011011010",
                      41 when "01010011011011",
                      41 when "01010011011100",
                      41 when "01010011011101",
                      41 when "01010011011110",
                      41 when "01010011011111",
                      41 when "01010011100000",
                      41 when "01010011100001",
                      41 when "01010011100010",
                      41 when "01010011100011",
                      41 when "01010011100100",
                      41 when "01010011100101",
                      41 when "01010011100110",
                      41 when "01010011100111",
                      41 when "01010011101000",
                      41 when "01010011101001",
                      41 when "01010011101010",
                      41 when "01010011101011",
                      41 when "01010011101100",
                      41 when "01010011101101",
                      41 when "01010011101110",
                      41 when "01010011101111",
                      41 when "01010011110000",
                      41 when "01010011110001",
                      41 when "01010011110010",
                      41 when "01010011110011",
                      41 when "01010011110100",
                      41 when "01010011110101",
                      41 when "01010011110110",
                      41 when "01010011110111",
                      41 when "01010011111000",
                      41 when "01010011111001",
                      41 when "01010011111010",
                      41 when "01010011111011",
                      41 when "01010011111100",
                      41 when "01010011111101",
                      41 when "01010011111110",
                      41 when "01010011111111",
                      41 when "01010100000000",
                      41 when "01010100000001",
                      41 when "01010100000010",
                      41 when "01010100000011",
                      41 when "01010100000100",
                      41 when "01010100000101",
                      41 when "01010100000110",
                      41 when "01010100000111",
                      41 when "01010100001000",
                      41 when "01010100001001",
                      41 when "01010100001010",
                      41 when "01010100001011",
                      41 when "01010100001100",
                      41 when "01010100001101",
                      41 when "01010100001110",
                      41 when "01010100001111",
                      41 when "01010100010000",
                      41 when "01010100010001",
                      41 when "01010100010010",
                      41 when "01010100010011",
                      41 when "01010100010100",
                      41 when "01010100010101",
                      41 when "01010100010110",
                      41 when "01010100010111",
                      41 when "01010100011000",
                      41 when "01010100011001",
                      41 when "01010100011010",
                      41 when "01010100011011",
                      41 when "01010100011100",
                      41 when "01010100011101",
                      41 when "01010100011110",
                      41 when "01010100011111",
                      41 when "01010100100000",
                      41 when "01010100100001",
                      41 when "01010100100010",
                      41 when "01010100100011",
                      41 when "01010100100100",
                      41 when "01010100100101",
                      41 when "01010100100110",
                      41 when "01010100100111",
                      41 when "01010100101000",
                      41 when "01010100101001",
                      41 when "01010100101010",
                      41 when "01010100101011",
                      41 when "01010100101100",
                      41 when "01010100101101",
                      41 when "01010100101110",
                      41 when "01010100101111",
                      41 when "01010100110000",
                      41 when "01010100110001",
                      40 when "01010100110010",
                      40 when "01010100110011",
                      40 when "01010100110100",
                      40 when "01010100110101",
                      40 when "01010100110110",
                      40 when "01010100110111",
                      40 when "01010100111000",
                      40 when "01010100111001",
                      40 when "01010100111010",
                      40 when "01010100111011",
                      40 when "01010100111100",
                      40 when "01010100111101",
                      40 when "01010100111110",
                      40 when "01010100111111",
                      40 when "01010101000000",
                      40 when "01010101000001",
                      40 when "01010101000010",
                      40 when "01010101000011",
                      40 when "01010101000100",
                      40 when "01010101000101",
                      40 when "01010101000110",
                      40 when "01010101000111",
                      40 when "01010101001000",
                      40 when "01010101001001",
                      40 when "01010101001010",
                      40 when "01010101001011",
                      40 when "01010101001100",
                      40 when "01010101001101",
                      40 when "01010101001110",
                      40 when "01010101001111",
                      40 when "01010101010000",
                      40 when "01010101010001",
                      40 when "01010101010010",
                      40 when "01010101010011",
                      40 when "01010101010100",
                      40 when "01010101010101",
                      40 when "01010101010110",
                      40 when "01010101010111",
                      40 when "01010101011000",
                      40 when "01010101011001",
                      40 when "01010101011010",
                      40 when "01010101011011",
                      40 when "01010101011100",
                      40 when "01010101011101",
                      40 when "01010101011110",
                      40 when "01010101011111",
                      40 when "01010101100000",
                      40 when "01010101100001",
                      40 when "01010101100010",
                      40 when "01010101100011",
                      40 when "01010101100100",
                      40 when "01010101100101",
                      40 when "01010101100110",
                      40 when "01010101100111",
                      40 when "01010101101000",
                      40 when "01010101101001",
                      40 when "01010101101010",
                      40 when "01010101101011",
                      40 when "01010101101100",
                      40 when "01010101101101",
                      40 when "01010101101110",
                      40 when "01010101101111",
                      40 when "01010101110000",
                      40 when "01010101110001",
                      40 when "01010101110010",
                      40 when "01010101110011",
                      40 when "01010101110100",
                      40 when "01010101110101",
                      40 when "01010101110110",
                      40 when "01010101110111",
                      40 when "01010101111000",
                      40 when "01010101111001",
                      40 when "01010101111010",
                      40 when "01010101111011",
                      40 when "01010101111100",
                      40 when "01010101111101",
                      40 when "01010101111110",
                      40 when "01010101111111",
                      40 when "01010110000000",
                      40 when "01010110000001",
                      40 when "01010110000010",
                      40 when "01010110000011",
                      40 when "01010110000100",
                      40 when "01010110000101",
                      40 when "01010110000110",
                      40 when "01010110000111",
                      40 when "01010110001000",
                      40 when "01010110001001",
                      40 when "01010110001010",
                      40 when "01010110001011",
                      40 when "01010110001100",
                      40 when "01010110001101",
                      40 when "01010110001110",
                      40 when "01010110001111",
                      40 when "01010110010000",
                      40 when "01010110010001",
                      40 when "01010110010010",
                      40 when "01010110010011",
                      40 when "01010110010100",
                      40 when "01010110010101",
                      40 when "01010110010110",
                      40 when "01010110010111",
                      40 when "01010110011000",
                      40 when "01010110011001",
                      40 when "01010110011010",
                      40 when "01010110011011",
                      40 when "01010110011100",
                      40 when "01010110011101",
                      40 when "01010110011110",
                      40 when "01010110011111",
                      40 when "01010110100000",
                      40 when "01010110100001",
                      40 when "01010110100010",
                      40 when "01010110100011",
                      40 when "01010110100100",
                      40 when "01010110100101",
                      40 when "01010110100110",
                      40 when "01010110100111",
                      40 when "01010110101000",
                      40 when "01010110101001",
                      40 when "01010110101010",
                      40 when "01010110101011",
                      40 when "01010110101100",
                      40 when "01010110101101",
                      40 when "01010110101110",
                      40 when "01010110101111",
                      40 when "01010110110000",
                      40 when "01010110110001",
                      40 when "01010110110010",
                      40 when "01010110110011",
                      40 when "01010110110100",
                      40 when "01010110110101",
                      40 when "01010110110110",
                      40 when "01010110110111",
                      40 when "01010110111000",
                      40 when "01010110111001",
                      40 when "01010110111010",
                      39 when "01010110111011",
                      39 when "01010110111100",
                      39 when "01010110111101",
                      39 when "01010110111110",
                      39 when "01010110111111",
                      39 when "01010111000000",
                      39 when "01010111000001",
                      39 when "01010111000010",
                      39 when "01010111000011",
                      39 when "01010111000100",
                      39 when "01010111000101",
                      39 when "01010111000110",
                      39 when "01010111000111",
                      39 when "01010111001000",
                      39 when "01010111001001",
                      39 when "01010111001010",
                      39 when "01010111001011",
                      39 when "01010111001100",
                      39 when "01010111001101",
                      39 when "01010111001110",
                      39 when "01010111001111",
                      39 when "01010111010000",
                      39 when "01010111010001",
                      39 when "01010111010010",
                      39 when "01010111010011",
                      39 when "01010111010100",
                      39 when "01010111010101",
                      39 when "01010111010110",
                      39 when "01010111010111",
                      39 when "01010111011000",
                      39 when "01010111011001",
                      39 when "01010111011010",
                      39 when "01010111011011",
                      39 when "01010111011100",
                      39 when "01010111011101",
                      39 when "01010111011110",
                      39 when "01010111011111",
                      39 when "01010111100000",
                      39 when "01010111100001",
                      39 when "01010111100010",
                      39 when "01010111100011",
                      39 when "01010111100100",
                      39 when "01010111100101",
                      39 when "01010111100110",
                      39 when "01010111100111",
                      39 when "01010111101000",
                      39 when "01010111101001",
                      39 when "01010111101010",
                      39 when "01010111101011",
                      39 when "01010111101100",
                      39 when "01010111101101",
                      39 when "01010111101110",
                      39 when "01010111101111",
                      39 when "01010111110000",
                      39 when "01010111110001",
                      39 when "01010111110010",
                      39 when "01010111110011",
                      39 when "01010111110100",
                      39 when "01010111110101",
                      39 when "01010111110110",
                      39 when "01010111110111",
                      39 when "01010111111000",
                      39 when "01010111111001",
                      39 when "01010111111010",
                      39 when "01010111111011",
                      39 when "01010111111100",
                      39 when "01010111111101",
                      39 when "01010111111110",
                      39 when "01010111111111",
                      39 when "01011000000000",
                      39 when "01011000000001",
                      39 when "01011000000010",
                      39 when "01011000000011",
                      39 when "01011000000100",
                      39 when "01011000000101",
                      39 when "01011000000110",
                      39 when "01011000000111",
                      39 when "01011000001000",
                      39 when "01011000001001",
                      39 when "01011000001010",
                      39 when "01011000001011",
                      39 when "01011000001100",
                      39 when "01011000001101",
                      39 when "01011000001110",
                      39 when "01011000001111",
                      39 when "01011000010000",
                      39 when "01011000010001",
                      39 when "01011000010010",
                      39 when "01011000010011",
                      39 when "01011000010100",
                      39 when "01011000010101",
                      39 when "01011000010110",
                      39 when "01011000010111",
                      39 when "01011000011000",
                      39 when "01011000011001",
                      39 when "01011000011010",
                      39 when "01011000011011",
                      39 when "01011000011100",
                      39 when "01011000011101",
                      39 when "01011000011110",
                      39 when "01011000011111",
                      39 when "01011000100000",
                      39 when "01011000100001",
                      39 when "01011000100010",
                      39 when "01011000100011",
                      39 when "01011000100100",
                      39 when "01011000100101",
                      39 when "01011000100110",
                      39 when "01011000100111",
                      39 when "01011000101000",
                      39 when "01011000101001",
                      39 when "01011000101010",
                      39 when "01011000101011",
                      39 when "01011000101100",
                      39 when "01011000101101",
                      39 when "01011000101110",
                      39 when "01011000101111",
                      39 when "01011000110000",
                      39 when "01011000110001",
                      39 when "01011000110010",
                      39 when "01011000110011",
                      39 when "01011000110100",
                      39 when "01011000110101",
                      39 when "01011000110110",
                      39 when "01011000110111",
                      39 when "01011000111000",
                      39 when "01011000111001",
                      39 when "01011000111010",
                      39 when "01011000111011",
                      39 when "01011000111100",
                      39 when "01011000111101",
                      39 when "01011000111110",
                      39 when "01011000111111",
                      39 when "01011001000000",
                      39 when "01011001000001",
                      39 when "01011001000010",
                      39 when "01011001000011",
                      39 when "01011001000100",
                      39 when "01011001000101",
                      39 when "01011001000110",
                      39 when "01011001000111",
                      39 when "01011001001000",
                      39 when "01011001001001",
                      39 when "01011001001010",
                      39 when "01011001001011",
                      38 when "01011001001100",
                      38 when "01011001001101",
                      38 when "01011001001110",
                      38 when "01011001001111",
                      38 when "01011001010000",
                      38 when "01011001010001",
                      38 when "01011001010010",
                      38 when "01011001010011",
                      38 when "01011001010100",
                      38 when "01011001010101",
                      38 when "01011001010110",
                      38 when "01011001010111",
                      38 when "01011001011000",
                      38 when "01011001011001",
                      38 when "01011001011010",
                      38 when "01011001011011",
                      38 when "01011001011100",
                      38 when "01011001011101",
                      38 when "01011001011110",
                      38 when "01011001011111",
                      38 when "01011001100000",
                      38 when "01011001100001",
                      38 when "01011001100010",
                      38 when "01011001100011",
                      38 when "01011001100100",
                      38 when "01011001100101",
                      38 when "01011001100110",
                      38 when "01011001100111",
                      38 when "01011001101000",
                      38 when "01011001101001",
                      38 when "01011001101010",
                      38 when "01011001101011",
                      38 when "01011001101100",
                      38 when "01011001101101",
                      38 when "01011001101110",
                      38 when "01011001101111",
                      38 when "01011001110000",
                      38 when "01011001110001",
                      38 when "01011001110010",
                      38 when "01011001110011",
                      38 when "01011001110100",
                      38 when "01011001110101",
                      38 when "01011001110110",
                      38 when "01011001110111",
                      38 when "01011001111000",
                      38 when "01011001111001",
                      38 when "01011001111010",
                      38 when "01011001111011",
                      38 when "01011001111100",
                      38 when "01011001111101",
                      38 when "01011001111110",
                      38 when "01011001111111",
                      38 when "01011010000000",
                      38 when "01011010000001",
                      38 when "01011010000010",
                      38 when "01011010000011",
                      38 when "01011010000100",
                      38 when "01011010000101",
                      38 when "01011010000110",
                      38 when "01011010000111",
                      38 when "01011010001000",
                      38 when "01011010001001",
                      38 when "01011010001010",
                      38 when "01011010001011",
                      38 when "01011010001100",
                      38 when "01011010001101",
                      38 when "01011010001110",
                      38 when "01011010001111",
                      38 when "01011010010000",
                      38 when "01011010010001",
                      38 when "01011010010010",
                      38 when "01011010010011",
                      38 when "01011010010100",
                      38 when "01011010010101",
                      38 when "01011010010110",
                      38 when "01011010010111",
                      38 when "01011010011000",
                      38 when "01011010011001",
                      38 when "01011010011010",
                      38 when "01011010011011",
                      38 when "01011010011100",
                      38 when "01011010011101",
                      38 when "01011010011110",
                      38 when "01011010011111",
                      38 when "01011010100000",
                      38 when "01011010100001",
                      38 when "01011010100010",
                      38 when "01011010100011",
                      38 when "01011010100100",
                      38 when "01011010100101",
                      38 when "01011010100110",
                      38 when "01011010100111",
                      38 when "01011010101000",
                      38 when "01011010101001",
                      38 when "01011010101010",
                      38 when "01011010101011",
                      38 when "01011010101100",
                      38 when "01011010101101",
                      38 when "01011010101110",
                      38 when "01011010101111",
                      38 when "01011010110000",
                      38 when "01011010110001",
                      38 when "01011010110010",
                      38 when "01011010110011",
                      38 when "01011010110100",
                      38 when "01011010110101",
                      38 when "01011010110110",
                      38 when "01011010110111",
                      38 when "01011010111000",
                      38 when "01011010111001",
                      38 when "01011010111010",
                      38 when "01011010111011",
                      38 when "01011010111100",
                      38 when "01011010111101",
                      38 when "01011010111110",
                      38 when "01011010111111",
                      38 when "01011011000000",
                      38 when "01011011000001",
                      38 when "01011011000010",
                      38 when "01011011000011",
                      38 when "01011011000100",
                      38 when "01011011000101",
                      38 when "01011011000110",
                      38 when "01011011000111",
                      38 when "01011011001000",
                      38 when "01011011001001",
                      38 when "01011011001010",
                      38 when "01011011001011",
                      38 when "01011011001100",
                      38 when "01011011001101",
                      38 when "01011011001110",
                      38 when "01011011001111",
                      38 when "01011011010000",
                      38 when "01011011010001",
                      38 when "01011011010010",
                      38 when "01011011010011",
                      38 when "01011011010100",
                      38 when "01011011010101",
                      38 when "01011011010110",
                      38 when "01011011010111",
                      38 when "01011011011000",
                      38 when "01011011011001",
                      38 when "01011011011010",
                      38 when "01011011011011",
                      38 when "01011011011100",
                      38 when "01011011011101",
                      38 when "01011011011110",
                      38 when "01011011011111",
                      38 when "01011011100000",
                      38 when "01011011100001",
                      38 when "01011011100010",
                      38 when "01011011100011",
                      37 when "01011011100100",
                      37 when "01011011100101",
                      37 when "01011011100110",
                      37 when "01011011100111",
                      37 when "01011011101000",
                      37 when "01011011101001",
                      37 when "01011011101010",
                      37 when "01011011101011",
                      37 when "01011011101100",
                      37 when "01011011101101",
                      37 when "01011011101110",
                      37 when "01011011101111",
                      37 when "01011011110000",
                      37 when "01011011110001",
                      37 when "01011011110010",
                      37 when "01011011110011",
                      37 when "01011011110100",
                      37 when "01011011110101",
                      37 when "01011011110110",
                      37 when "01011011110111",
                      37 when "01011011111000",
                      37 when "01011011111001",
                      37 when "01011011111010",
                      37 when "01011011111011",
                      37 when "01011011111100",
                      37 when "01011011111101",
                      37 when "01011011111110",
                      37 when "01011011111111",
                      37 when "01011100000000",
                      37 when "01011100000001",
                      37 when "01011100000010",
                      37 when "01011100000011",
                      37 when "01011100000100",
                      37 when "01011100000101",
                      37 when "01011100000110",
                      37 when "01011100000111",
                      37 when "01011100001000",
                      37 when "01011100001001",
                      37 when "01011100001010",
                      37 when "01011100001011",
                      37 when "01011100001100",
                      37 when "01011100001101",
                      37 when "01011100001110",
                      37 when "01011100001111",
                      37 when "01011100010000",
                      37 when "01011100010001",
                      37 when "01011100010010",
                      37 when "01011100010011",
                      37 when "01011100010100",
                      37 when "01011100010101",
                      37 when "01011100010110",
                      37 when "01011100010111",
                      37 when "01011100011000",
                      37 when "01011100011001",
                      37 when "01011100011010",
                      37 when "01011100011011",
                      37 when "01011100011100",
                      37 when "01011100011101",
                      37 when "01011100011110",
                      37 when "01011100011111",
                      37 when "01011100100000",
                      37 when "01011100100001",
                      37 when "01011100100010",
                      37 when "01011100100011",
                      37 when "01011100100100",
                      37 when "01011100100101",
                      37 when "01011100100110",
                      37 when "01011100100111",
                      37 when "01011100101000",
                      37 when "01011100101001",
                      37 when "01011100101010",
                      37 when "01011100101011",
                      37 when "01011100101100",
                      37 when "01011100101101",
                      37 when "01011100101110",
                      37 when "01011100101111",
                      37 when "01011100110000",
                      37 when "01011100110001",
                      37 when "01011100110010",
                      37 when "01011100110011",
                      37 when "01011100110100",
                      37 when "01011100110101",
                      37 when "01011100110110",
                      37 when "01011100110111",
                      37 when "01011100111000",
                      37 when "01011100111001",
                      37 when "01011100111010",
                      37 when "01011100111011",
                      37 when "01011100111100",
                      37 when "01011100111101",
                      37 when "01011100111110",
                      37 when "01011100111111",
                      37 when "01011101000000",
                      37 when "01011101000001",
                      37 when "01011101000010",
                      37 when "01011101000011",
                      37 when "01011101000100",
                      37 when "01011101000101",
                      37 when "01011101000110",
                      37 when "01011101000111",
                      37 when "01011101001000",
                      37 when "01011101001001",
                      37 when "01011101001010",
                      37 when "01011101001011",
                      37 when "01011101001100",
                      37 when "01011101001101",
                      37 when "01011101001110",
                      37 when "01011101001111",
                      37 when "01011101010000",
                      37 when "01011101010001",
                      37 when "01011101010010",
                      37 when "01011101010011",
                      37 when "01011101010100",
                      37 when "01011101010101",
                      37 when "01011101010110",
                      37 when "01011101010111",
                      37 when "01011101011000",
                      37 when "01011101011001",
                      37 when "01011101011010",
                      37 when "01011101011011",
                      37 when "01011101011100",
                      37 when "01011101011101",
                      37 when "01011101011110",
                      37 when "01011101011111",
                      37 when "01011101100000",
                      37 when "01011101100001",
                      37 when "01011101100010",
                      37 when "01011101100011",
                      37 when "01011101100100",
                      37 when "01011101100101",
                      37 when "01011101100110",
                      37 when "01011101100111",
                      37 when "01011101101000",
                      37 when "01011101101001",
                      37 when "01011101101010",
                      37 when "01011101101011",
                      37 when "01011101101100",
                      37 when "01011101101101",
                      37 when "01011101101110",
                      37 when "01011101101111",
                      37 when "01011101110000",
                      37 when "01011101110001",
                      37 when "01011101110010",
                      37 when "01011101110011",
                      37 when "01011101110100",
                      37 when "01011101110101",
                      37 when "01011101110110",
                      37 when "01011101110111",
                      37 when "01011101111000",
                      37 when "01011101111001",
                      37 when "01011101111010",
                      37 when "01011101111011",
                      37 when "01011101111100",
                      37 when "01011101111101",
                      37 when "01011101111110",
                      37 when "01011101111111",
                      37 when "01011110000000",
                      37 when "01011110000001",
                      37 when "01011110000010",
                      37 when "01011110000011",
                      36 when "01011110000100",
                      36 when "01011110000101",
                      36 when "01011110000110",
                      36 when "01011110000111",
                      36 when "01011110001000",
                      36 when "01011110001001",
                      36 when "01011110001010",
                      36 when "01011110001011",
                      36 when "01011110001100",
                      36 when "01011110001101",
                      36 when "01011110001110",
                      36 when "01011110001111",
                      36 when "01011110010000",
                      36 when "01011110010001",
                      36 when "01011110010010",
                      36 when "01011110010011",
                      36 when "01011110010100",
                      36 when "01011110010101",
                      36 when "01011110010110",
                      36 when "01011110010111",
                      36 when "01011110011000",
                      36 when "01011110011001",
                      36 when "01011110011010",
                      36 when "01011110011011",
                      36 when "01011110011100",
                      36 when "01011110011101",
                      36 when "01011110011110",
                      36 when "01011110011111",
                      36 when "01011110100000",
                      36 when "01011110100001",
                      36 when "01011110100010",
                      36 when "01011110100011",
                      36 when "01011110100100",
                      36 when "01011110100101",
                      36 when "01011110100110",
                      36 when "01011110100111",
                      36 when "01011110101000",
                      36 when "01011110101001",
                      36 when "01011110101010",
                      36 when "01011110101011",
                      36 when "01011110101100",
                      36 when "01011110101101",
                      36 when "01011110101110",
                      36 when "01011110101111",
                      36 when "01011110110000",
                      36 when "01011110110001",
                      36 when "01011110110010",
                      36 when "01011110110011",
                      36 when "01011110110100",
                      36 when "01011110110101",
                      36 when "01011110110110",
                      36 when "01011110110111",
                      36 when "01011110111000",
                      36 when "01011110111001",
                      36 when "01011110111010",
                      36 when "01011110111011",
                      36 when "01011110111100",
                      36 when "01011110111101",
                      36 when "01011110111110",
                      36 when "01011110111111",
                      36 when "01011111000000",
                      36 when "01011111000001",
                      36 when "01011111000010",
                      36 when "01011111000011",
                      36 when "01011111000100",
                      36 when "01011111000101",
                      36 when "01011111000110",
                      36 when "01011111000111",
                      36 when "01011111001000",
                      36 when "01011111001001",
                      36 when "01011111001010",
                      36 when "01011111001011",
                      36 when "01011111001100",
                      36 when "01011111001101",
                      36 when "01011111001110",
                      36 when "01011111001111",
                      36 when "01011111010000",
                      36 when "01011111010001",
                      36 when "01011111010010",
                      36 when "01011111010011",
                      36 when "01011111010100",
                      36 when "01011111010101",
                      36 when "01011111010110",
                      36 when "01011111010111",
                      36 when "01011111011000",
                      36 when "01011111011001",
                      36 when "01011111011010",
                      36 when "01011111011011",
                      36 when "01011111011100",
                      36 when "01011111011101",
                      36 when "01011111011110",
                      36 when "01011111011111",
                      36 when "01011111100000",
                      36 when "01011111100001",
                      36 when "01011111100010",
                      36 when "01011111100011",
                      36 when "01011111100100",
                      36 when "01011111100101",
                      36 when "01011111100110",
                      36 when "01011111100111",
                      36 when "01011111101000",
                      36 when "01011111101001",
                      36 when "01011111101010",
                      36 when "01011111101011",
                      36 when "01011111101100",
                      36 when "01011111101101",
                      36 when "01011111101110",
                      36 when "01011111101111",
                      36 when "01011111110000",
                      36 when "01011111110001",
                      36 when "01011111110010",
                      36 when "01011111110011",
                      36 when "01011111110100",
                      36 when "01011111110101",
                      36 when "01011111110110",
                      36 when "01011111110111",
                      36 when "01011111111000",
                      36 when "01011111111001",
                      36 when "01011111111010",
                      36 when "01011111111011",
                      36 when "01011111111100",
                      36 when "01011111111101",
                      36 when "01011111111110",
                      36 when "01011111111111",
                      36 when "01100000000000",
                      36 when "01100000000001",
                      36 when "01100000000010",
                      36 when "01100000000011",
                      36 when "01100000000100",
                      36 when "01100000000101",
                      36 when "01100000000110",
                      36 when "01100000000111",
                      36 when "01100000001000",
                      36 when "01100000001001",
                      36 when "01100000001010",
                      36 when "01100000001011",
                      36 when "01100000001100",
                      36 when "01100000001101",
                      36 when "01100000001110",
                      36 when "01100000001111",
                      36 when "01100000010000",
                      36 when "01100000010001",
                      36 when "01100000010010",
                      36 when "01100000010011",
                      36 when "01100000010100",
                      36 when "01100000010101",
                      36 when "01100000010110",
                      36 when "01100000010111",
                      36 when "01100000011000",
                      36 when "01100000011001",
                      36 when "01100000011010",
                      36 when "01100000011011",
                      36 when "01100000011100",
                      36 when "01100000011101",
                      36 when "01100000011110",
                      36 when "01100000011111",
                      36 when "01100000100000",
                      36 when "01100000100001",
                      36 when "01100000100010",
                      36 when "01100000100011",
                      36 when "01100000100100",
                      36 when "01100000100101",
                      36 when "01100000100110",
                      36 when "01100000100111",
                      36 when "01100000101000",
                      36 when "01100000101001",
                      36 when "01100000101010",
                      36 when "01100000101011",
                      36 when "01100000101100",
                      36 when "01100000101101",
                      35 when "01100000101110",
                      35 when "01100000101111",
                      35 when "01100000110000",
                      35 when "01100000110001",
                      35 when "01100000110010",
                      35 when "01100000110011",
                      35 when "01100000110100",
                      35 when "01100000110101",
                      35 when "01100000110110",
                      35 when "01100000110111",
                      35 when "01100000111000",
                      35 when "01100000111001",
                      35 when "01100000111010",
                      35 when "01100000111011",
                      35 when "01100000111100",
                      35 when "01100000111101",
                      35 when "01100000111110",
                      35 when "01100000111111",
                      35 when "01100001000000",
                      35 when "01100001000001",
                      35 when "01100001000010",
                      35 when "01100001000011",
                      35 when "01100001000100",
                      35 when "01100001000101",
                      35 when "01100001000110",
                      35 when "01100001000111",
                      35 when "01100001001000",
                      35 when "01100001001001",
                      35 when "01100001001010",
                      35 when "01100001001011",
                      35 when "01100001001100",
                      35 when "01100001001101",
                      35 when "01100001001110",
                      35 when "01100001001111",
                      35 when "01100001010000",
                      35 when "01100001010001",
                      35 when "01100001010010",
                      35 when "01100001010011",
                      35 when "01100001010100",
                      35 when "01100001010101",
                      35 when "01100001010110",
                      35 when "01100001010111",
                      35 when "01100001011000",
                      35 when "01100001011001",
                      35 when "01100001011010",
                      35 when "01100001011011",
                      35 when "01100001011100",
                      35 when "01100001011101",
                      35 when "01100001011110",
                      35 when "01100001011111",
                      35 when "01100001100000",
                      35 when "01100001100001",
                      35 when "01100001100010",
                      35 when "01100001100011",
                      35 when "01100001100100",
                      35 when "01100001100101",
                      35 when "01100001100110",
                      35 when "01100001100111",
                      35 when "01100001101000",
                      35 when "01100001101001",
                      35 when "01100001101010",
                      35 when "01100001101011",
                      35 when "01100001101100",
                      35 when "01100001101101",
                      35 when "01100001101110",
                      35 when "01100001101111",
                      35 when "01100001110000",
                      35 when "01100001110001",
                      35 when "01100001110010",
                      35 when "01100001110011",
                      35 when "01100001110100",
                      35 when "01100001110101",
                      35 when "01100001110110",
                      35 when "01100001110111",
                      35 when "01100001111000",
                      35 when "01100001111001",
                      35 when "01100001111010",
                      35 when "01100001111011",
                      35 when "01100001111100",
                      35 when "01100001111101",
                      35 when "01100001111110",
                      35 when "01100001111111",
                      35 when "01100010000000",
                      35 when "01100010000001",
                      35 when "01100010000010",
                      35 when "01100010000011",
                      35 when "01100010000100",
                      35 when "01100010000101",
                      35 when "01100010000110",
                      35 when "01100010000111",
                      35 when "01100010001000",
                      35 when "01100010001001",
                      35 when "01100010001010",
                      35 when "01100010001011",
                      35 when "01100010001100",
                      35 when "01100010001101",
                      35 when "01100010001110",
                      35 when "01100010001111",
                      35 when "01100010010000",
                      35 when "01100010010001",
                      35 when "01100010010010",
                      35 when "01100010010011",
                      35 when "01100010010100",
                      35 when "01100010010101",
                      35 when "01100010010110",
                      35 when "01100010010111",
                      35 when "01100010011000",
                      35 when "01100010011001",
                      35 when "01100010011010",
                      35 when "01100010011011",
                      35 when "01100010011100",
                      35 when "01100010011101",
                      35 when "01100010011110",
                      35 when "01100010011111",
                      35 when "01100010100000",
                      35 when "01100010100001",
                      35 when "01100010100010",
                      35 when "01100010100011",
                      35 when "01100010100100",
                      35 when "01100010100101",
                      35 when "01100010100110",
                      35 when "01100010100111",
                      35 when "01100010101000",
                      35 when "01100010101001",
                      35 when "01100010101010",
                      35 when "01100010101011",
                      35 when "01100010101100",
                      35 when "01100010101101",
                      35 when "01100010101110",
                      35 when "01100010101111",
                      35 when "01100010110000",
                      35 when "01100010110001",
                      35 when "01100010110010",
                      35 when "01100010110011",
                      35 when "01100010110100",
                      35 when "01100010110101",
                      35 when "01100010110110",
                      35 when "01100010110111",
                      35 when "01100010111000",
                      35 when "01100010111001",
                      35 when "01100010111010",
                      35 when "01100010111011",
                      35 when "01100010111100",
                      35 when "01100010111101",
                      35 when "01100010111110",
                      35 when "01100010111111",
                      35 when "01100011000000",
                      35 when "01100011000001",
                      35 when "01100011000010",
                      35 when "01100011000011",
                      35 when "01100011000100",
                      35 when "01100011000101",
                      35 when "01100011000110",
                      35 when "01100011000111",
                      35 when "01100011001000",
                      35 when "01100011001001",
                      35 when "01100011001010",
                      35 when "01100011001011",
                      35 when "01100011001100",
                      35 when "01100011001101",
                      35 when "01100011001110",
                      35 when "01100011001111",
                      35 when "01100011010000",
                      35 when "01100011010001",
                      35 when "01100011010010",
                      35 when "01100011010011",
                      35 when "01100011010100",
                      35 when "01100011010101",
                      35 when "01100011010110",
                      35 when "01100011010111",
                      35 when "01100011011000",
                      35 when "01100011011001",
                      35 when "01100011011010",
                      35 when "01100011011011",
                      35 when "01100011011100",
                      35 when "01100011011101",
                      35 when "01100011011110",
                      35 when "01100011011111",
                      35 when "01100011100000",
                      34 when "01100011100001",
                      34 when "01100011100010",
                      34 when "01100011100011",
                      34 when "01100011100100",
                      34 when "01100011100101",
                      34 when "01100011100110",
                      34 when "01100011100111",
                      34 when "01100011101000",
                      34 when "01100011101001",
                      34 when "01100011101010",
                      34 when "01100011101011",
                      34 when "01100011101100",
                      34 when "01100011101101",
                      34 when "01100011101110",
                      34 when "01100011101111",
                      34 when "01100011110000",
                      34 when "01100011110001",
                      34 when "01100011110010",
                      34 when "01100011110011",
                      34 when "01100011110100",
                      34 when "01100011110101",
                      34 when "01100011110110",
                      34 when "01100011110111",
                      34 when "01100011111000",
                      34 when "01100011111001",
                      34 when "01100011111010",
                      34 when "01100011111011",
                      34 when "01100011111100",
                      34 when "01100011111101",
                      34 when "01100011111110",
                      34 when "01100011111111",
                      34 when "01100100000000",
                      34 when "01100100000001",
                      34 when "01100100000010",
                      34 when "01100100000011",
                      34 when "01100100000100",
                      34 when "01100100000101",
                      34 when "01100100000110",
                      34 when "01100100000111",
                      34 when "01100100001000",
                      34 when "01100100001001",
                      34 when "01100100001010",
                      34 when "01100100001011",
                      34 when "01100100001100",
                      34 when "01100100001101",
                      34 when "01100100001110",
                      34 when "01100100001111",
                      34 when "01100100010000",
                      34 when "01100100010001",
                      34 when "01100100010010",
                      34 when "01100100010011",
                      34 when "01100100010100",
                      34 when "01100100010101",
                      34 when "01100100010110",
                      34 when "01100100010111",
                      34 when "01100100011000",
                      34 when "01100100011001",
                      34 when "01100100011010",
                      34 when "01100100011011",
                      34 when "01100100011100",
                      34 when "01100100011101",
                      34 when "01100100011110",
                      34 when "01100100011111",
                      34 when "01100100100000",
                      34 when "01100100100001",
                      34 when "01100100100010",
                      34 when "01100100100011",
                      34 when "01100100100100",
                      34 when "01100100100101",
                      34 when "01100100100110",
                      34 when "01100100100111",
                      34 when "01100100101000",
                      34 when "01100100101001",
                      34 when "01100100101010",
                      34 when "01100100101011",
                      34 when "01100100101100",
                      34 when "01100100101101",
                      34 when "01100100101110",
                      34 when "01100100101111",
                      34 when "01100100110000",
                      34 when "01100100110001",
                      34 when "01100100110010",
                      34 when "01100100110011",
                      34 when "01100100110100",
                      34 when "01100100110101",
                      34 when "01100100110110",
                      34 when "01100100110111",
                      34 when "01100100111000",
                      34 when "01100100111001",
                      34 when "01100100111010",
                      34 when "01100100111011",
                      34 when "01100100111100",
                      34 when "01100100111101",
                      34 when "01100100111110",
                      34 when "01100100111111",
                      34 when "01100101000000",
                      34 when "01100101000001",
                      34 when "01100101000010",
                      34 when "01100101000011",
                      34 when "01100101000100",
                      34 when "01100101000101",
                      34 when "01100101000110",
                      34 when "01100101000111",
                      34 when "01100101001000",
                      34 when "01100101001001",
                      34 when "01100101001010",
                      34 when "01100101001011",
                      34 when "01100101001100",
                      34 when "01100101001101",
                      34 when "01100101001110",
                      34 when "01100101001111",
                      34 when "01100101010000",
                      34 when "01100101010001",
                      34 when "01100101010010",
                      34 when "01100101010011",
                      34 when "01100101010100",
                      34 when "01100101010101",
                      34 when "01100101010110",
                      34 when "01100101010111",
                      34 when "01100101011000",
                      34 when "01100101011001",
                      34 when "01100101011010",
                      34 when "01100101011011",
                      34 when "01100101011100",
                      34 when "01100101011101",
                      34 when "01100101011110",
                      34 when "01100101011111",
                      34 when "01100101100000",
                      34 when "01100101100001",
                      34 when "01100101100010",
                      34 when "01100101100011",
                      34 when "01100101100100",
                      34 when "01100101100101",
                      34 when "01100101100110",
                      34 when "01100101100111",
                      34 when "01100101101000",
                      34 when "01100101101001",
                      34 when "01100101101010",
                      34 when "01100101101011",
                      34 when "01100101101100",
                      34 when "01100101101101",
                      34 when "01100101101110",
                      34 when "01100101101111",
                      34 when "01100101110000",
                      34 when "01100101110001",
                      34 when "01100101110010",
                      34 when "01100101110011",
                      34 when "01100101110100",
                      34 when "01100101110101",
                      34 when "01100101110110",
                      34 when "01100101110111",
                      34 when "01100101111000",
                      34 when "01100101111001",
                      34 when "01100101111010",
                      34 when "01100101111011",
                      34 when "01100101111100",
                      34 when "01100101111101",
                      34 when "01100101111110",
                      34 when "01100101111111",
                      34 when "01100110000000",
                      34 when "01100110000001",
                      34 when "01100110000010",
                      34 when "01100110000011",
                      34 when "01100110000100",
                      34 when "01100110000101",
                      34 when "01100110000110",
                      34 when "01100110000111",
                      34 when "01100110001000",
                      34 when "01100110001001",
                      34 when "01100110001010",
                      34 when "01100110001011",
                      34 when "01100110001100",
                      34 when "01100110001101",
                      34 when "01100110001110",
                      34 when "01100110001111",
                      34 when "01100110010000",
                      34 when "01100110010001",
                      34 when "01100110010010",
                      34 when "01100110010011",
                      34 when "01100110010100",
                      34 when "01100110010101",
                      34 when "01100110010110",
                      34 when "01100110010111",
                      34 when "01100110011000",
                      34 when "01100110011001",
                      34 when "01100110011010",
                      34 when "01100110011011",
                      34 when "01100110011100",
                      34 when "01100110011101",
                      34 when "01100110011110",
                      34 when "01100110011111",
                      33 when "01100110100000",
                      33 when "01100110100001",
                      33 when "01100110100010",
                      33 when "01100110100011",
                      33 when "01100110100100",
                      33 when "01100110100101",
                      33 when "01100110100110",
                      33 when "01100110100111",
                      33 when "01100110101000",
                      33 when "01100110101001",
                      33 when "01100110101010",
                      33 when "01100110101011",
                      33 when "01100110101100",
                      33 when "01100110101101",
                      33 when "01100110101110",
                      33 when "01100110101111",
                      33 when "01100110110000",
                      33 when "01100110110001",
                      33 when "01100110110010",
                      33 when "01100110110011",
                      33 when "01100110110100",
                      33 when "01100110110101",
                      33 when "01100110110110",
                      33 when "01100110110111",
                      33 when "01100110111000",
                      33 when "01100110111001",
                      33 when "01100110111010",
                      33 when "01100110111011",
                      33 when "01100110111100",
                      33 when "01100110111101",
                      33 when "01100110111110",
                      33 when "01100110111111",
                      33 when "01100111000000",
                      33 when "01100111000001",
                      33 when "01100111000010",
                      33 when "01100111000011",
                      33 when "01100111000100",
                      33 when "01100111000101",
                      33 when "01100111000110",
                      33 when "01100111000111",
                      33 when "01100111001000",
                      33 when "01100111001001",
                      33 when "01100111001010",
                      33 when "01100111001011",
                      33 when "01100111001100",
                      33 when "01100111001101",
                      33 when "01100111001110",
                      33 when "01100111001111",
                      33 when "01100111010000",
                      33 when "01100111010001",
                      33 when "01100111010010",
                      33 when "01100111010011",
                      33 when "01100111010100",
                      33 when "01100111010101",
                      33 when "01100111010110",
                      33 when "01100111010111",
                      33 when "01100111011000",
                      33 when "01100111011001",
                      33 when "01100111011010",
                      33 when "01100111011011",
                      33 when "01100111011100",
                      33 when "01100111011101",
                      33 when "01100111011110",
                      33 when "01100111011111",
                      33 when "01100111100000",
                      33 when "01100111100001",
                      33 when "01100111100010",
                      33 when "01100111100011",
                      33 when "01100111100100",
                      33 when "01100111100101",
                      33 when "01100111100110",
                      33 when "01100111100111",
                      33 when "01100111101000",
                      33 when "01100111101001",
                      33 when "01100111101010",
                      33 when "01100111101011",
                      33 when "01100111101100",
                      33 when "01100111101101",
                      33 when "01100111101110",
                      33 when "01100111101111",
                      33 when "01100111110000",
                      33 when "01100111110001",
                      33 when "01100111110010",
                      33 when "01100111110011",
                      33 when "01100111110100",
                      33 when "01100111110101",
                      33 when "01100111110110",
                      33 when "01100111110111",
                      33 when "01100111111000",
                      33 when "01100111111001",
                      33 when "01100111111010",
                      33 when "01100111111011",
                      33 when "01100111111100",
                      33 when "01100111111101",
                      33 when "01100111111110",
                      33 when "01100111111111",
                      33 when "01101000000000",
                      33 when "01101000000001",
                      33 when "01101000000010",
                      33 when "01101000000011",
                      33 when "01101000000100",
                      33 when "01101000000101",
                      33 when "01101000000110",
                      33 when "01101000000111",
                      33 when "01101000001000",
                      33 when "01101000001001",
                      33 when "01101000001010",
                      33 when "01101000001011",
                      33 when "01101000001100",
                      33 when "01101000001101",
                      33 when "01101000001110",
                      33 when "01101000001111",
                      33 when "01101000010000",
                      33 when "01101000010001",
                      33 when "01101000010010",
                      33 when "01101000010011",
                      33 when "01101000010100",
                      33 when "01101000010101",
                      33 when "01101000010110",
                      33 when "01101000010111",
                      33 when "01101000011000",
                      33 when "01101000011001",
                      33 when "01101000011010",
                      33 when "01101000011011",
                      33 when "01101000011100",
                      33 when "01101000011101",
                      33 when "01101000011110",
                      33 when "01101000011111",
                      33 when "01101000100000",
                      33 when "01101000100001",
                      33 when "01101000100010",
                      33 when "01101000100011",
                      33 when "01101000100100",
                      33 when "01101000100101",
                      33 when "01101000100110",
                      33 when "01101000100111",
                      33 when "01101000101000",
                      33 when "01101000101001",
                      33 when "01101000101010",
                      33 when "01101000101011",
                      33 when "01101000101100",
                      33 when "01101000101101",
                      33 when "01101000101110",
                      33 when "01101000101111",
                      33 when "01101000110000",
                      33 when "01101000110001",
                      33 when "01101000110010",
                      33 when "01101000110011",
                      33 when "01101000110100",
                      33 when "01101000110101",
                      33 when "01101000110110",
                      33 when "01101000110111",
                      33 when "01101000111000",
                      33 when "01101000111001",
                      33 when "01101000111010",
                      33 when "01101000111011",
                      33 when "01101000111100",
                      33 when "01101000111101",
                      33 when "01101000111110",
                      33 when "01101000111111",
                      33 when "01101001000000",
                      33 when "01101001000001",
                      33 when "01101001000010",
                      33 when "01101001000011",
                      33 when "01101001000100",
                      33 when "01101001000101",
                      33 when "01101001000110",
                      33 when "01101001000111",
                      33 when "01101001001000",
                      33 when "01101001001001",
                      33 when "01101001001010",
                      33 when "01101001001011",
                      33 when "01101001001100",
                      33 when "01101001001101",
                      33 when "01101001001110",
                      33 when "01101001001111",
                      33 when "01101001010000",
                      33 when "01101001010001",
                      33 when "01101001010010",
                      33 when "01101001010011",
                      33 when "01101001010100",
                      33 when "01101001010101",
                      33 when "01101001010110",
                      33 when "01101001010111",
                      33 when "01101001011000",
                      33 when "01101001011001",
                      33 when "01101001011010",
                      33 when "01101001011011",
                      33 when "01101001011100",
                      33 when "01101001011101",
                      33 when "01101001011110",
                      33 when "01101001011111",
                      33 when "01101001100000",
                      33 when "01101001100001",
                      33 when "01101001100010",
                      33 when "01101001100011",
                      33 when "01101001100100",
                      33 when "01101001100101",
                      33 when "01101001100110",
                      33 when "01101001100111",
                      33 when "01101001101000",
                      32 when "01101001101001",
                      32 when "01101001101010",
                      32 when "01101001101011",
                      32 when "01101001101100",
                      32 when "01101001101101",
                      32 when "01101001101110",
                      32 when "01101001101111",
                      32 when "01101001110000",
                      32 when "01101001110001",
                      32 when "01101001110010",
                      32 when "01101001110011",
                      32 when "01101001110100",
                      32 when "01101001110101",
                      32 when "01101001110110",
                      32 when "01101001110111",
                      32 when "01101001111000",
                      32 when "01101001111001",
                      32 when "01101001111010",
                      32 when "01101001111011",
                      32 when "01101001111100",
                      32 when "01101001111101",
                      32 when "01101001111110",
                      32 when "01101001111111",
                      32 when "01101010000000",
                      32 when "01101010000001",
                      32 when "01101010000010",
                      32 when "01101010000011",
                      32 when "01101010000100",
                      32 when "01101010000101",
                      32 when "01101010000110",
                      32 when "01101010000111",
                      32 when "01101010001000",
                      32 when "01101010001001",
                      32 when "01101010001010",
                      32 when "01101010001011",
                      32 when "01101010001100",
                      32 when "01101010001101",
                      32 when "01101010001110",
                      32 when "01101010001111",
                      32 when "01101010010000",
                      32 when "01101010010001",
                      32 when "01101010010010",
                      32 when "01101010010011",
                      32 when "01101010010100",
                      32 when "01101010010101",
                      32 when "01101010010110",
                      32 when "01101010010111",
                      32 when "01101010011000",
                      32 when "01101010011001",
                      32 when "01101010011010",
                      32 when "01101010011011",
                      32 when "01101010011100",
                      32 when "01101010011101",
                      32 when "01101010011110",
                      32 when "01101010011111",
                      32 when "01101010100000",
                      32 when "01101010100001",
                      32 when "01101010100010",
                      32 when "01101010100011",
                      32 when "01101010100100",
                      32 when "01101010100101",
                      32 when "01101010100110",
                      32 when "01101010100111",
                      32 when "01101010101000",
                      32 when "01101010101001",
                      32 when "01101010101010",
                      32 when "01101010101011",
                      32 when "01101010101100",
                      32 when "01101010101101",
                      32 when "01101010101110",
                      32 when "01101010101111",
                      32 when "01101010110000",
                      32 when "01101010110001",
                      32 when "01101010110010",
                      32 when "01101010110011",
                      32 when "01101010110100",
                      32 when "01101010110101",
                      32 when "01101010110110",
                      32 when "01101010110111",
                      32 when "01101010111000",
                      32 when "01101010111001",
                      32 when "01101010111010",
                      32 when "01101010111011",
                      32 when "01101010111100",
                      32 when "01101010111101",
                      32 when "01101010111110",
                      32 when "01101010111111",
                      32 when "01101011000000",
                      32 when "01101011000001",
                      32 when "01101011000010",
                      32 when "01101011000011",
                      32 when "01101011000100",
                      32 when "01101011000101",
                      32 when "01101011000110",
                      32 when "01101011000111",
                      32 when "01101011001000",
                      32 when "01101011001001",
                      32 when "01101011001010",
                      32 when "01101011001011",
                      32 when "01101011001100",
                      32 when "01101011001101",
                      32 when "01101011001110",
                      32 when "01101011001111",
                      32 when "01101011010000",
                      32 when "01101011010001",
                      32 when "01101011010010",
                      32 when "01101011010011",
                      32 when "01101011010100",
                      32 when "01101011010101",
                      32 when "01101011010110",
                      32 when "01101011010111",
                      32 when "01101011011000",
                      32 when "01101011011001",
                      32 when "01101011011010",
                      32 when "01101011011011",
                      32 when "01101011011100",
                      32 when "01101011011101",
                      32 when "01101011011110",
                      32 when "01101011011111",
                      32 when "01101011100000",
                      32 when "01101011100001",
                      32 when "01101011100010",
                      32 when "01101011100011",
                      32 when "01101011100100",
                      32 when "01101011100101",
                      32 when "01101011100110",
                      32 when "01101011100111",
                      32 when "01101011101000",
                      32 when "01101011101001",
                      32 when "01101011101010",
                      32 when "01101011101011",
                      32 when "01101011101100",
                      32 when "01101011101101",
                      32 when "01101011101110",
                      32 when "01101011101111",
                      32 when "01101011110000",
                      32 when "01101011110001",
                      32 when "01101011110010",
                      32 when "01101011110011",
                      32 when "01101011110100",
                      32 when "01101011110101",
                      32 when "01101011110110",
                      32 when "01101011110111",
                      32 when "01101011111000",
                      32 when "01101011111001",
                      32 when "01101011111010",
                      32 when "01101011111011",
                      32 when "01101011111100",
                      32 when "01101011111101",
                      32 when "01101011111110",
                      32 when "01101011111111",
                      32 when "01101100000000",
                      32 when "01101100000001",
                      32 when "01101100000010",
                      32 when "01101100000011",
                      32 when "01101100000100",
                      32 when "01101100000101",
                      32 when "01101100000110",
                      32 when "01101100000111",
                      32 when "01101100001000",
                      32 when "01101100001001",
                      32 when "01101100001010",
                      32 when "01101100001011",
                      32 when "01101100001100",
                      32 when "01101100001101",
                      32 when "01101100001110",
                      32 when "01101100001111",
                      32 when "01101100010000",
                      32 when "01101100010001",
                      32 when "01101100010010",
                      32 when "01101100010011",
                      32 when "01101100010100",
                      32 when "01101100010101",
                      32 when "01101100010110",
                      32 when "01101100010111",
                      32 when "01101100011000",
                      32 when "01101100011001",
                      32 when "01101100011010",
                      32 when "01101100011011",
                      32 when "01101100011100",
                      32 when "01101100011101",
                      32 when "01101100011110",
                      32 when "01101100011111",
                      32 when "01101100100000",
                      32 when "01101100100001",
                      32 when "01101100100010",
                      32 when "01101100100011",
                      32 when "01101100100100",
                      32 when "01101100100101",
                      32 when "01101100100110",
                      32 when "01101100100111",
                      32 when "01101100101000",
                      32 when "01101100101001",
                      32 when "01101100101010",
                      32 when "01101100101011",
                      32 when "01101100101100",
                      32 when "01101100101101",
                      32 when "01101100101110",
                      32 when "01101100101111",
                      32 when "01101100110000",
                      32 when "01101100110001",
                      32 when "01101100110010",
                      32 when "01101100110011",
                      32 when "01101100110100",
                      32 when "01101100110101",
                      32 when "01101100110110",
                      32 when "01101100110111",
                      32 when "01101100111000",
                      32 when "01101100111001",
                      32 when "01101100111010",
                      32 when "01101100111011",
                      32 when "01101100111100",
                      32 when "01101100111101",
                      32 when "01101100111110",
                      32 when "01101100111111",
                      31 when "01101101000000",
                      31 when "01101101000001",
                      31 when "01101101000010",
                      31 when "01101101000011",
                      31 when "01101101000100",
                      31 when "01101101000101",
                      31 when "01101101000110",
                      31 when "01101101000111",
                      31 when "01101101001000",
                      31 when "01101101001001",
                      31 when "01101101001010",
                      31 when "01101101001011",
                      31 when "01101101001100",
                      31 when "01101101001101",
                      31 when "01101101001110",
                      31 when "01101101001111",
                      31 when "01101101010000",
                      31 when "01101101010001",
                      31 when "01101101010010",
                      31 when "01101101010011",
                      31 when "01101101010100",
                      31 when "01101101010101",
                      31 when "01101101010110",
                      31 when "01101101010111",
                      31 when "01101101011000",
                      31 when "01101101011001",
                      31 when "01101101011010",
                      31 when "01101101011011",
                      31 when "01101101011100",
                      31 when "01101101011101",
                      31 when "01101101011110",
                      31 when "01101101011111",
                      31 when "01101101100000",
                      31 when "01101101100001",
                      31 when "01101101100010",
                      31 when "01101101100011",
                      31 when "01101101100100",
                      31 when "01101101100101",
                      31 when "01101101100110",
                      31 when "01101101100111",
                      31 when "01101101101000",
                      31 when "01101101101001",
                      31 when "01101101101010",
                      31 when "01101101101011",
                      31 when "01101101101100",
                      31 when "01101101101101",
                      31 when "01101101101110",
                      31 when "01101101101111",
                      31 when "01101101110000",
                      31 when "01101101110001",
                      31 when "01101101110010",
                      31 when "01101101110011",
                      31 when "01101101110100",
                      31 when "01101101110101",
                      31 when "01101101110110",
                      31 when "01101101110111",
                      31 when "01101101111000",
                      31 when "01101101111001",
                      31 when "01101101111010",
                      31 when "01101101111011",
                      31 when "01101101111100",
                      31 when "01101101111101",
                      31 when "01101101111110",
                      31 when "01101101111111",
                      31 when "01101110000000",
                      31 when "01101110000001",
                      31 when "01101110000010",
                      31 when "01101110000011",
                      31 when "01101110000100",
                      31 when "01101110000101",
                      31 when "01101110000110",
                      31 when "01101110000111",
                      31 when "01101110001000",
                      31 when "01101110001001",
                      31 when "01101110001010",
                      31 when "01101110001011",
                      31 when "01101110001100",
                      31 when "01101110001101",
                      31 when "01101110001110",
                      31 when "01101110001111",
                      31 when "01101110010000",
                      31 when "01101110010001",
                      31 when "01101110010010",
                      31 when "01101110010011",
                      31 when "01101110010100",
                      31 when "01101110010101",
                      31 when "01101110010110",
                      31 when "01101110010111",
                      31 when "01101110011000",
                      31 when "01101110011001",
                      31 when "01101110011010",
                      31 when "01101110011011",
                      31 when "01101110011100",
                      31 when "01101110011101",
                      31 when "01101110011110",
                      31 when "01101110011111",
                      31 when "01101110100000",
                      31 when "01101110100001",
                      31 when "01101110100010",
                      31 when "01101110100011",
                      31 when "01101110100100",
                      31 when "01101110100101",
                      31 when "01101110100110",
                      31 when "01101110100111",
                      31 when "01101110101000",
                      31 when "01101110101001",
                      31 when "01101110101010",
                      31 when "01101110101011",
                      31 when "01101110101100",
                      31 when "01101110101101",
                      31 when "01101110101110",
                      31 when "01101110101111",
                      31 when "01101110110000",
                      31 when "01101110110001",
                      31 when "01101110110010",
                      31 when "01101110110011",
                      31 when "01101110110100",
                      31 when "01101110110101",
                      31 when "01101110110110",
                      31 when "01101110110111",
                      31 when "01101110111000",
                      31 when "01101110111001",
                      31 when "01101110111010",
                      31 when "01101110111011",
                      31 when "01101110111100",
                      31 when "01101110111101",
                      31 when "01101110111110",
                      31 when "01101110111111",
                      31 when "01101111000000",
                      31 when "01101111000001",
                      31 when "01101111000010",
                      31 when "01101111000011",
                      31 when "01101111000100",
                      31 when "01101111000101",
                      31 when "01101111000110",
                      31 when "01101111000111",
                      31 when "01101111001000",
                      31 when "01101111001001",
                      31 when "01101111001010",
                      31 when "01101111001011",
                      31 when "01101111001100",
                      31 when "01101111001101",
                      31 when "01101111001110",
                      31 when "01101111001111",
                      31 when "01101111010000",
                      31 when "01101111010001",
                      31 when "01101111010010",
                      31 when "01101111010011",
                      31 when "01101111010100",
                      31 when "01101111010101",
                      31 when "01101111010110",
                      31 when "01101111010111",
                      31 when "01101111011000",
                      31 when "01101111011001",
                      31 when "01101111011010",
                      31 when "01101111011011",
                      31 when "01101111011100",
                      31 when "01101111011101",
                      31 when "01101111011110",
                      31 when "01101111011111",
                      31 when "01101111100000",
                      31 when "01101111100001",
                      31 when "01101111100010",
                      31 when "01101111100011",
                      31 when "01101111100100",
                      31 when "01101111100101",
                      31 when "01101111100110",
                      31 when "01101111100111",
                      31 when "01101111101000",
                      31 when "01101111101001",
                      31 when "01101111101010",
                      31 when "01101111101011",
                      31 when "01101111101100",
                      31 when "01101111101101",
                      31 when "01101111101110",
                      31 when "01101111101111",
                      31 when "01101111110000",
                      31 when "01101111110001",
                      31 when "01101111110010",
                      31 when "01101111110011",
                      31 when "01101111110100",
                      31 when "01101111110101",
                      31 when "01101111110110",
                      31 when "01101111110111",
                      31 when "01101111111000",
                      31 when "01101111111001",
                      31 when "01101111111010",
                      31 when "01101111111011",
                      31 when "01101111111100",
                      31 when "01101111111101",
                      31 when "01101111111110",
                      31 when "01101111111111",
                      31 when "01110000000000",
                      31 when "01110000000001",
                      31 when "01110000000010",
                      31 when "01110000000011",
                      31 when "01110000000100",
                      31 when "01110000000101",
                      31 when "01110000000110",
                      31 when "01110000000111",
                      31 when "01110000001000",
                      31 when "01110000001001",
                      31 when "01110000001010",
                      31 when "01110000001011",
                      31 when "01110000001100",
                      31 when "01110000001101",
                      31 when "01110000001110",
                      31 when "01110000001111",
                      31 when "01110000010000",
                      31 when "01110000010001",
                      31 when "01110000010010",
                      31 when "01110000010011",
                      31 when "01110000010100",
                      31 when "01110000010101",
                      31 when "01110000010110",
                      31 when "01110000010111",
                      31 when "01110000011000",
                      31 when "01110000011001",
                      31 when "01110000011010",
                      31 when "01110000011011",
                      31 when "01110000011100",
                      31 when "01110000011101",
                      31 when "01110000011110",
                      31 when "01110000011111",
                      31 when "01110000100000",
                      31 when "01110000100001",
                      31 when "01110000100010",
                      31 when "01110000100011",
                      31 when "01110000100100",
                      30 when "01110000100101",
                      30 when "01110000100110",
                      30 when "01110000100111",
                      30 when "01110000101000",
                      30 when "01110000101001",
                      30 when "01110000101010",
                      30 when "01110000101011",
                      30 when "01110000101100",
                      30 when "01110000101101",
                      30 when "01110000101110",
                      30 when "01110000101111",
                      30 when "01110000110000",
                      30 when "01110000110001",
                      30 when "01110000110010",
                      30 when "01110000110011",
                      30 when "01110000110100",
                      30 when "01110000110101",
                      30 when "01110000110110",
                      30 when "01110000110111",
                      30 when "01110000111000",
                      30 when "01110000111001",
                      30 when "01110000111010",
                      30 when "01110000111011",
                      30 when "01110000111100",
                      30 when "01110000111101",
                      30 when "01110000111110",
                      30 when "01110000111111",
                      30 when "01110001000000",
                      30 when "01110001000001",
                      30 when "01110001000010",
                      30 when "01110001000011",
                      30 when "01110001000100",
                      30 when "01110001000101",
                      30 when "01110001000110",
                      30 when "01110001000111",
                      30 when "01110001001000",
                      30 when "01110001001001",
                      30 when "01110001001010",
                      30 when "01110001001011",
                      30 when "01110001001100",
                      30 when "01110001001101",
                      30 when "01110001001110",
                      30 when "01110001001111",
                      30 when "01110001010000",
                      30 when "01110001010001",
                      30 when "01110001010010",
                      30 when "01110001010011",
                      30 when "01110001010100",
                      30 when "01110001010101",
                      30 when "01110001010110",
                      30 when "01110001010111",
                      30 when "01110001011000",
                      30 when "01110001011001",
                      30 when "01110001011010",
                      30 when "01110001011011",
                      30 when "01110001011100",
                      30 when "01110001011101",
                      30 when "01110001011110",
                      30 when "01110001011111",
                      30 when "01110001100000",
                      30 when "01110001100001",
                      30 when "01110001100010",
                      30 when "01110001100011",
                      30 when "01110001100100",
                      30 when "01110001100101",
                      30 when "01110001100110",
                      30 when "01110001100111",
                      30 when "01110001101000",
                      30 when "01110001101001",
                      30 when "01110001101010",
                      30 when "01110001101011",
                      30 when "01110001101100",
                      30 when "01110001101101",
                      30 when "01110001101110",
                      30 when "01110001101111",
                      30 when "01110001110000",
                      30 when "01110001110001",
                      30 when "01110001110010",
                      30 when "01110001110011",
                      30 when "01110001110100",
                      30 when "01110001110101",
                      30 when "01110001110110",
                      30 when "01110001110111",
                      30 when "01110001111000",
                      30 when "01110001111001",
                      30 when "01110001111010",
                      30 when "01110001111011",
                      30 when "01110001111100",
                      30 when "01110001111101",
                      30 when "01110001111110",
                      30 when "01110001111111",
                      30 when "01110010000000",
                      30 when "01110010000001",
                      30 when "01110010000010",
                      30 when "01110010000011",
                      30 when "01110010000100",
                      30 when "01110010000101",
                      30 when "01110010000110",
                      30 when "01110010000111",
                      30 when "01110010001000",
                      30 when "01110010001001",
                      30 when "01110010001010",
                      30 when "01110010001011",
                      30 when "01110010001100",
                      30 when "01110010001101",
                      30 when "01110010001110",
                      30 when "01110010001111",
                      30 when "01110010010000",
                      30 when "01110010010001",
                      30 when "01110010010010",
                      30 when "01110010010011",
                      30 when "01110010010100",
                      30 when "01110010010101",
                      30 when "01110010010110",
                      30 when "01110010010111",
                      30 when "01110010011000",
                      30 when "01110010011001",
                      30 when "01110010011010",
                      30 when "01110010011011",
                      30 when "01110010011100",
                      30 when "01110010011101",
                      30 when "01110010011110",
                      30 when "01110010011111",
                      30 when "01110010100000",
                      30 when "01110010100001",
                      30 when "01110010100010",
                      30 when "01110010100011",
                      30 when "01110010100100",
                      30 when "01110010100101",
                      30 when "01110010100110",
                      30 when "01110010100111",
                      30 when "01110010101000",
                      30 when "01110010101001",
                      30 when "01110010101010",
                      30 when "01110010101011",
                      30 when "01110010101100",
                      30 when "01110010101101",
                      30 when "01110010101110",
                      30 when "01110010101111",
                      30 when "01110010110000",
                      30 when "01110010110001",
                      30 when "01110010110010",
                      30 when "01110010110011",
                      30 when "01110010110100",
                      30 when "01110010110101",
                      30 when "01110010110110",
                      30 when "01110010110111",
                      30 when "01110010111000",
                      30 when "01110010111001",
                      30 when "01110010111010",
                      30 when "01110010111011",
                      30 when "01110010111100",
                      30 when "01110010111101",
                      30 when "01110010111110",
                      30 when "01110010111111",
                      30 when "01110011000000",
                      30 when "01110011000001",
                      30 when "01110011000010",
                      30 when "01110011000011",
                      30 when "01110011000100",
                      30 when "01110011000101",
                      30 when "01110011000110",
                      30 when "01110011000111",
                      30 when "01110011001000",
                      30 when "01110011001001",
                      30 when "01110011001010",
                      30 when "01110011001011",
                      30 when "01110011001100",
                      30 when "01110011001101",
                      30 when "01110011001110",
                      30 when "01110011001111",
                      30 when "01110011010000",
                      30 when "01110011010001",
                      30 when "01110011010010",
                      30 when "01110011010011",
                      30 when "01110011010100",
                      30 when "01110011010101",
                      30 when "01110011010110",
                      30 when "01110011010111",
                      30 when "01110011011000",
                      30 when "01110011011001",
                      30 when "01110011011010",
                      30 when "01110011011011",
                      30 when "01110011011100",
                      30 when "01110011011101",
                      30 when "01110011011110",
                      30 when "01110011011111",
                      30 when "01110011100000",
                      30 when "01110011100001",
                      30 when "01110011100010",
                      30 when "01110011100011",
                      30 when "01110011100100",
                      30 when "01110011100101",
                      30 when "01110011100110",
                      30 when "01110011100111",
                      30 when "01110011101000",
                      30 when "01110011101001",
                      30 when "01110011101010",
                      30 when "01110011101011",
                      30 when "01110011101100",
                      30 when "01110011101101",
                      30 when "01110011101110",
                      30 when "01110011101111",
                      30 when "01110011110000",
                      30 when "01110011110001",
                      30 when "01110011110010",
                      30 when "01110011110011",
                      30 when "01110011110100",
                      30 when "01110011110101",
                      30 when "01110011110110",
                      30 when "01110011110111",
                      30 when "01110011111000",
                      30 when "01110011111001",
                      30 when "01110011111010",
                      30 when "01110011111011",
                      30 when "01110011111100",
                      30 when "01110011111101",
                      30 when "01110011111110",
                      30 when "01110011111111",
                      30 when "01110100000000",
                      30 when "01110100000001",
                      30 when "01110100000010",
                      30 when "01110100000011",
                      30 when "01110100000100",
                      30 when "01110100000101",
                      30 when "01110100000110",
                      30 when "01110100000111",
                      30 when "01110100001000",
                      30 when "01110100001001",
                      30 when "01110100001010",
                      30 when "01110100001011",
                      30 when "01110100001100",
                      30 when "01110100001101",
                      30 when "01110100001110",
                      30 when "01110100001111",
                      30 when "01110100010000",
                      30 when "01110100010001",
                      30 when "01110100010010",
                      30 when "01110100010011",
                      30 when "01110100010100",
                      30 when "01110100010101",
                      30 when "01110100010110",
                      30 when "01110100010111",
                      30 when "01110100011000",
                      29 when "01110100011001",
                      29 when "01110100011010",
                      29 when "01110100011011",
                      29 when "01110100011100",
                      29 when "01110100011101",
                      29 when "01110100011110",
                      29 when "01110100011111",
                      29 when "01110100100000",
                      29 when "01110100100001",
                      29 when "01110100100010",
                      29 when "01110100100011",
                      29 when "01110100100100",
                      29 when "01110100100101",
                      29 when "01110100100110",
                      29 when "01110100100111",
                      29 when "01110100101000",
                      29 when "01110100101001",
                      29 when "01110100101010",
                      29 when "01110100101011",
                      29 when "01110100101100",
                      29 when "01110100101101",
                      29 when "01110100101110",
                      29 when "01110100101111",
                      29 when "01110100110000",
                      29 when "01110100110001",
                      29 when "01110100110010",
                      29 when "01110100110011",
                      29 when "01110100110100",
                      29 when "01110100110101",
                      29 when "01110100110110",
                      29 when "01110100110111",
                      29 when "01110100111000",
                      29 when "01110100111001",
                      29 when "01110100111010",
                      29 when "01110100111011",
                      29 when "01110100111100",
                      29 when "01110100111101",
                      29 when "01110100111110",
                      29 when "01110100111111",
                      29 when "01110101000000",
                      29 when "01110101000001",
                      29 when "01110101000010",
                      29 when "01110101000011",
                      29 when "01110101000100",
                      29 when "01110101000101",
                      29 when "01110101000110",
                      29 when "01110101000111",
                      29 when "01110101001000",
                      29 when "01110101001001",
                      29 when "01110101001010",
                      29 when "01110101001011",
                      29 when "01110101001100",
                      29 when "01110101001101",
                      29 when "01110101001110",
                      29 when "01110101001111",
                      29 when "01110101010000",
                      29 when "01110101010001",
                      29 when "01110101010010",
                      29 when "01110101010011",
                      29 when "01110101010100",
                      29 when "01110101010101",
                      29 when "01110101010110",
                      29 when "01110101010111",
                      29 when "01110101011000",
                      29 when "01110101011001",
                      29 when "01110101011010",
                      29 when "01110101011011",
                      29 when "01110101011100",
                      29 when "01110101011101",
                      29 when "01110101011110",
                      29 when "01110101011111",
                      29 when "01110101100000",
                      29 when "01110101100001",
                      29 when "01110101100010",
                      29 when "01110101100011",
                      29 when "01110101100100",
                      29 when "01110101100101",
                      29 when "01110101100110",
                      29 when "01110101100111",
                      29 when "01110101101000",
                      29 when "01110101101001",
                      29 when "01110101101010",
                      29 when "01110101101011",
                      29 when "01110101101100",
                      29 when "01110101101101",
                      29 when "01110101101110",
                      29 when "01110101101111",
                      29 when "01110101110000",
                      29 when "01110101110001",
                      29 when "01110101110010",
                      29 when "01110101110011",
                      29 when "01110101110100",
                      29 when "01110101110101",
                      29 when "01110101110110",
                      29 when "01110101110111",
                      29 when "01110101111000",
                      29 when "01110101111001",
                      29 when "01110101111010",
                      29 when "01110101111011",
                      29 when "01110101111100",
                      29 when "01110101111101",
                      29 when "01110101111110",
                      29 when "01110101111111",
                      29 when "01110110000000",
                      29 when "01110110000001",
                      29 when "01110110000010",
                      29 when "01110110000011",
                      29 when "01110110000100",
                      29 when "01110110000101",
                      29 when "01110110000110",
                      29 when "01110110000111",
                      29 when "01110110001000",
                      29 when "01110110001001",
                      29 when "01110110001010",
                      29 when "01110110001011",
                      29 when "01110110001100",
                      29 when "01110110001101",
                      29 when "01110110001110",
                      29 when "01110110001111",
                      29 when "01110110010000",
                      29 when "01110110010001",
                      29 when "01110110010010",
                      29 when "01110110010011",
                      29 when "01110110010100",
                      29 when "01110110010101",
                      29 when "01110110010110",
                      29 when "01110110010111",
                      29 when "01110110011000",
                      29 when "01110110011001",
                      29 when "01110110011010",
                      29 when "01110110011011",
                      29 when "01110110011100",
                      29 when "01110110011101",
                      29 when "01110110011110",
                      29 when "01110110011111",
                      29 when "01110110100000",
                      29 when "01110110100001",
                      29 when "01110110100010",
                      29 when "01110110100011",
                      29 when "01110110100100",
                      29 when "01110110100101",
                      29 when "01110110100110",
                      29 when "01110110100111",
                      29 when "01110110101000",
                      29 when "01110110101001",
                      29 when "01110110101010",
                      29 when "01110110101011",
                      29 when "01110110101100",
                      29 when "01110110101101",
                      29 when "01110110101110",
                      29 when "01110110101111",
                      29 when "01110110110000",
                      29 when "01110110110001",
                      29 when "01110110110010",
                      29 when "01110110110011",
                      29 when "01110110110100",
                      29 when "01110110110101",
                      29 when "01110110110110",
                      29 when "01110110110111",
                      29 when "01110110111000",
                      29 when "01110110111001",
                      29 when "01110110111010",
                      29 when "01110110111011",
                      29 when "01110110111100",
                      29 when "01110110111101",
                      29 when "01110110111110",
                      29 when "01110110111111",
                      29 when "01110111000000",
                      29 when "01110111000001",
                      29 when "01110111000010",
                      29 when "01110111000011",
                      29 when "01110111000100",
                      29 when "01110111000101",
                      29 when "01110111000110",
                      29 when "01110111000111",
                      29 when "01110111001000",
                      29 when "01110111001001",
                      29 when "01110111001010",
                      29 when "01110111001011",
                      29 when "01110111001100",
                      29 when "01110111001101",
                      29 when "01110111001110",
                      29 when "01110111001111",
                      29 when "01110111010000",
                      29 when "01110111010001",
                      29 when "01110111010010",
                      29 when "01110111010011",
                      29 when "01110111010100",
                      29 when "01110111010101",
                      29 when "01110111010110",
                      29 when "01110111010111",
                      29 when "01110111011000",
                      29 when "01110111011001",
                      29 when "01110111011010",
                      29 when "01110111011011",
                      29 when "01110111011100",
                      29 when "01110111011101",
                      29 when "01110111011110",
                      29 when "01110111011111",
                      29 when "01110111100000",
                      29 when "01110111100001",
                      29 when "01110111100010",
                      29 when "01110111100011",
                      29 when "01110111100100",
                      29 when "01110111100101",
                      29 when "01110111100110",
                      29 when "01110111100111",
                      29 when "01110111101000",
                      29 when "01110111101001",
                      29 when "01110111101010",
                      29 when "01110111101011",
                      29 when "01110111101100",
                      29 when "01110111101101",
                      29 when "01110111101110",
                      29 when "01110111101111",
                      29 when "01110111110000",
                      29 when "01110111110001",
                      29 when "01110111110010",
                      29 when "01110111110011",
                      29 when "01110111110100",
                      29 when "01110111110101",
                      29 when "01110111110110",
                      29 when "01110111110111",
                      29 when "01110111111000",
                      29 when "01110111111001",
                      29 when "01110111111010",
                      29 when "01110111111011",
                      29 when "01110111111100",
                      29 when "01110111111101",
                      29 when "01110111111110",
                      29 when "01110111111111",
                      29 when "01111000000000",
                      29 when "01111000000001",
                      29 when "01111000000010",
                      29 when "01111000000011",
                      29 when "01111000000100",
                      29 when "01111000000101",
                      29 when "01111000000110",
                      29 when "01111000000111",
                      29 when "01111000001000",
                      29 when "01111000001001",
                      29 when "01111000001010",
                      29 when "01111000001011",
                      29 when "01111000001100",
                      29 when "01111000001101",
                      29 when "01111000001110",
                      29 when "01111000001111",
                      29 when "01111000010000",
                      29 when "01111000010001",
                      29 when "01111000010010",
                      29 when "01111000010011",
                      29 when "01111000010100",
                      29 when "01111000010101",
                      29 when "01111000010110",
                      29 when "01111000010111",
                      29 when "01111000011000",
                      29 when "01111000011001",
                      29 when "01111000011010",
                      29 when "01111000011011",
                      29 when "01111000011100",
                      29 when "01111000011101",
                      28 when "01111000011110",
                      28 when "01111000011111",
                      28 when "01111000100000",
                      28 when "01111000100001",
                      28 when "01111000100010",
                      28 when "01111000100011",
                      28 when "01111000100100",
                      28 when "01111000100101",
                      28 when "01111000100110",
                      28 when "01111000100111",
                      28 when "01111000101000",
                      28 when "01111000101001",
                      28 when "01111000101010",
                      28 when "01111000101011",
                      28 when "01111000101100",
                      28 when "01111000101101",
                      28 when "01111000101110",
                      28 when "01111000101111",
                      28 when "01111000110000",
                      28 when "01111000110001",
                      28 when "01111000110010",
                      28 when "01111000110011",
                      28 when "01111000110100",
                      28 when "01111000110101",
                      28 when "01111000110110",
                      28 when "01111000110111",
                      28 when "01111000111000",
                      28 when "01111000111001",
                      28 when "01111000111010",
                      28 when "01111000111011",
                      28 when "01111000111100",
                      28 when "01111000111101",
                      28 when "01111000111110",
                      28 when "01111000111111",
                      28 when "01111001000000",
                      28 when "01111001000001",
                      28 when "01111001000010",
                      28 when "01111001000011",
                      28 when "01111001000100",
                      28 when "01111001000101",
                      28 when "01111001000110",
                      28 when "01111001000111",
                      28 when "01111001001000",
                      28 when "01111001001001",
                      28 when "01111001001010",
                      28 when "01111001001011",
                      28 when "01111001001100",
                      28 when "01111001001101",
                      28 when "01111001001110",
                      28 when "01111001001111",
                      28 when "01111001010000",
                      28 when "01111001010001",
                      28 when "01111001010010",
                      28 when "01111001010011",
                      28 when "01111001010100",
                      28 when "01111001010101",
                      28 when "01111001010110",
                      28 when "01111001010111",
                      28 when "01111001011000",
                      28 when "01111001011001",
                      28 when "01111001011010",
                      28 when "01111001011011",
                      28 when "01111001011100",
                      28 when "01111001011101",
                      28 when "01111001011110",
                      28 when "01111001011111",
                      28 when "01111001100000",
                      28 when "01111001100001",
                      28 when "01111001100010",
                      28 when "01111001100011",
                      28 when "01111001100100",
                      28 when "01111001100101",
                      28 when "01111001100110",
                      28 when "01111001100111",
                      28 when "01111001101000",
                      28 when "01111001101001",
                      28 when "01111001101010",
                      28 when "01111001101011",
                      28 when "01111001101100",
                      28 when "01111001101101",
                      28 when "01111001101110",
                      28 when "01111001101111",
                      28 when "01111001110000",
                      28 when "01111001110001",
                      28 when "01111001110010",
                      28 when "01111001110011",
                      28 when "01111001110100",
                      28 when "01111001110101",
                      28 when "01111001110110",
                      28 when "01111001110111",
                      28 when "01111001111000",
                      28 when "01111001111001",
                      28 when "01111001111010",
                      28 when "01111001111011",
                      28 when "01111001111100",
                      28 when "01111001111101",
                      28 when "01111001111110",
                      28 when "01111001111111",
                      28 when "01111010000000",
                      28 when "01111010000001",
                      28 when "01111010000010",
                      28 when "01111010000011",
                      28 when "01111010000100",
                      28 when "01111010000101",
                      28 when "01111010000110",
                      28 when "01111010000111",
                      28 when "01111010001000",
                      28 when "01111010001001",
                      28 when "01111010001010",
                      28 when "01111010001011",
                      28 when "01111010001100",
                      28 when "01111010001101",
                      28 when "01111010001110",
                      28 when "01111010001111",
                      28 when "01111010010000",
                      28 when "01111010010001",
                      28 when "01111010010010",
                      28 when "01111010010011",
                      28 when "01111010010100",
                      28 when "01111010010101",
                      28 when "01111010010110",
                      28 when "01111010010111",
                      28 when "01111010011000",
                      28 when "01111010011001",
                      28 when "01111010011010",
                      28 when "01111010011011",
                      28 when "01111010011100",
                      28 when "01111010011101",
                      28 when "01111010011110",
                      28 when "01111010011111",
                      28 when "01111010100000",
                      28 when "01111010100001",
                      28 when "01111010100010",
                      28 when "01111010100011",
                      28 when "01111010100100",
                      28 when "01111010100101",
                      28 when "01111010100110",
                      28 when "01111010100111",
                      28 when "01111010101000",
                      28 when "01111010101001",
                      28 when "01111010101010",
                      28 when "01111010101011",
                      28 when "01111010101100",
                      28 when "01111010101101",
                      28 when "01111010101110",
                      28 when "01111010101111",
                      28 when "01111010110000",
                      28 when "01111010110001",
                      28 when "01111010110010",
                      28 when "01111010110011",
                      28 when "01111010110100",
                      28 when "01111010110101",
                      28 when "01111010110110",
                      28 when "01111010110111",
                      28 when "01111010111000",
                      28 when "01111010111001",
                      28 when "01111010111010",
                      28 when "01111010111011",
                      28 when "01111010111100",
                      28 when "01111010111101",
                      28 when "01111010111110",
                      28 when "01111010111111",
                      28 when "01111011000000",
                      28 when "01111011000001",
                      28 when "01111011000010",
                      28 when "01111011000011",
                      28 when "01111011000100",
                      28 when "01111011000101",
                      28 when "01111011000110",
                      28 when "01111011000111",
                      28 when "01111011001000",
                      28 when "01111011001001",
                      28 when "01111011001010",
                      28 when "01111011001011",
                      28 when "01111011001100",
                      28 when "01111011001101",
                      28 when "01111011001110",
                      28 when "01111011001111",
                      28 when "01111011010000",
                      28 when "01111011010001",
                      28 when "01111011010010",
                      28 when "01111011010011",
                      28 when "01111011010100",
                      28 when "01111011010101",
                      28 when "01111011010110",
                      28 when "01111011010111",
                      28 when "01111011011000",
                      28 when "01111011011001",
                      28 when "01111011011010",
                      28 when "01111011011011",
                      28 when "01111011011100",
                      28 when "01111011011101",
                      28 when "01111011011110",
                      28 when "01111011011111",
                      28 when "01111011100000",
                      28 when "01111011100001",
                      28 when "01111011100010",
                      28 when "01111011100011",
                      28 when "01111011100100",
                      28 when "01111011100101",
                      28 when "01111011100110",
                      28 when "01111011100111",
                      28 when "01111011101000",
                      28 when "01111011101001",
                      28 when "01111011101010",
                      28 when "01111011101011",
                      28 when "01111011101100",
                      28 when "01111011101101",
                      28 when "01111011101110",
                      28 when "01111011101111",
                      28 when "01111011110000",
                      28 when "01111011110001",
                      28 when "01111011110010",
                      28 when "01111011110011",
                      28 when "01111011110100",
                      28 when "01111011110101",
                      28 when "01111011110110",
                      28 when "01111011110111",
                      28 when "01111011111000",
                      28 when "01111011111001",
                      28 when "01111011111010",
                      28 when "01111011111011",
                      28 when "01111011111100",
                      28 when "01111011111101",
                      28 when "01111011111110",
                      28 when "01111011111111",
                      28 when "01111100000000",
                      28 when "01111100000001",
                      28 when "01111100000010",
                      28 when "01111100000011",
                      28 when "01111100000100",
                      28 when "01111100000101",
                      28 when "01111100000110",
                      28 when "01111100000111",
                      28 when "01111100001000",
                      28 when "01111100001001",
                      28 when "01111100001010",
                      28 when "01111100001011",
                      28 when "01111100001100",
                      28 when "01111100001101",
                      28 when "01111100001110",
                      28 when "01111100001111",
                      28 when "01111100010000",
                      28 when "01111100010001",
                      28 when "01111100010010",
                      28 when "01111100010011",
                      28 when "01111100010100",
                      28 when "01111100010101",
                      28 when "01111100010110",
                      28 when "01111100010111",
                      28 when "01111100011000",
                      28 when "01111100011001",
                      28 when "01111100011010",
                      28 when "01111100011011",
                      28 when "01111100011100",
                      28 when "01111100011101",
                      28 when "01111100011110",
                      28 when "01111100011111",
                      28 when "01111100100000",
                      28 when "01111100100001",
                      28 when "01111100100010",
                      28 when "01111100100011",
                      28 when "01111100100100",
                      28 when "01111100100101",
                      28 when "01111100100110",
                      28 when "01111100100111",
                      28 when "01111100101000",
                      28 when "01111100101001",
                      28 when "01111100101010",
                      28 when "01111100101011",
                      28 when "01111100101100",
                      28 when "01111100101101",
                      28 when "01111100101110",
                      28 when "01111100101111",
                      28 when "01111100110000",
                      28 when "01111100110001",
                      28 when "01111100110010",
                      28 when "01111100110011",
                      28 when "01111100110100",
                      28 when "01111100110101",
                      28 when "01111100110110",
                      27 when "01111100110111",
                      27 when "01111100111000",
                      27 when "01111100111001",
                      27 when "01111100111010",
                      27 when "01111100111011",
                      27 when "01111100111100",
                      27 when "01111100111101",
                      27 when "01111100111110",
                      27 when "01111100111111",
                      27 when "01111101000000",
                      27 when "01111101000001",
                      27 when "01111101000010",
                      27 when "01111101000011",
                      27 when "01111101000100",
                      27 when "01111101000101",
                      27 when "01111101000110",
                      27 when "01111101000111",
                      27 when "01111101001000",
                      27 when "01111101001001",
                      27 when "01111101001010",
                      27 when "01111101001011",
                      27 when "01111101001100",
                      27 when "01111101001101",
                      27 when "01111101001110",
                      27 when "01111101001111",
                      27 when "01111101010000",
                      27 when "01111101010001",
                      27 when "01111101010010",
                      27 when "01111101010011",
                      27 when "01111101010100",
                      27 when "01111101010101",
                      27 when "01111101010110",
                      27 when "01111101010111",
                      27 when "01111101011000",
                      27 when "01111101011001",
                      27 when "01111101011010",
                      27 when "01111101011011",
                      27 when "01111101011100",
                      27 when "01111101011101",
                      27 when "01111101011110",
                      27 when "01111101011111",
                      27 when "01111101100000",
                      27 when "01111101100001",
                      27 when "01111101100010",
                      27 when "01111101100011",
                      27 when "01111101100100",
                      27 when "01111101100101",
                      27 when "01111101100110",
                      27 when "01111101100111",
                      27 when "01111101101000",
                      27 when "01111101101001",
                      27 when "01111101101010",
                      27 when "01111101101011",
                      27 when "01111101101100",
                      27 when "01111101101101",
                      27 when "01111101101110",
                      27 when "01111101101111",
                      27 when "01111101110000",
                      27 when "01111101110001",
                      27 when "01111101110010",
                      27 when "01111101110011",
                      27 when "01111101110100",
                      27 when "01111101110101",
                      27 when "01111101110110",
                      27 when "01111101110111",
                      27 when "01111101111000",
                      27 when "01111101111001",
                      27 when "01111101111010",
                      27 when "01111101111011",
                      27 when "01111101111100",
                      27 when "01111101111101",
                      27 when "01111101111110",
                      27 when "01111101111111",
                      27 when "01111110000000",
                      27 when "01111110000001",
                      27 when "01111110000010",
                      27 when "01111110000011",
                      27 when "01111110000100",
                      27 when "01111110000101",
                      27 when "01111110000110",
                      27 when "01111110000111",
                      27 when "01111110001000",
                      27 when "01111110001001",
                      27 when "01111110001010",
                      27 when "01111110001011",
                      27 when "01111110001100",
                      27 when "01111110001101",
                      27 when "01111110001110",
                      27 when "01111110001111",
                      27 when "01111110010000",
                      27 when "01111110010001",
                      27 when "01111110010010",
                      27 when "01111110010011",
                      27 when "01111110010100",
                      27 when "01111110010101",
                      27 when "01111110010110",
                      27 when "01111110010111",
                      27 when "01111110011000",
                      27 when "01111110011001",
                      27 when "01111110011010",
                      27 when "01111110011011",
                      27 when "01111110011100",
                      27 when "01111110011101",
                      27 when "01111110011110",
                      27 when "01111110011111",
                      27 when "01111110100000",
                      27 when "01111110100001",
                      27 when "01111110100010",
                      27 when "01111110100011",
                      27 when "01111110100100",
                      27 when "01111110100101",
                      27 when "01111110100110",
                      27 when "01111110100111",
                      27 when "01111110101000",
                      27 when "01111110101001",
                      27 when "01111110101010",
                      27 when "01111110101011",
                      27 when "01111110101100",
                      27 when "01111110101101",
                      27 when "01111110101110",
                      27 when "01111110101111",
                      27 when "01111110110000",
                      27 when "01111110110001",
                      27 when "01111110110010",
                      27 when "01111110110011",
                      27 when "01111110110100",
                      27 when "01111110110101",
                      27 when "01111110110110",
                      27 when "01111110110111",
                      27 when "01111110111000",
                      27 when "01111110111001",
                      27 when "01111110111010",
                      27 when "01111110111011",
                      27 when "01111110111100",
                      27 when "01111110111101",
                      27 when "01111110111110",
                      27 when "01111110111111",
                      27 when "01111111000000",
                      27 when "01111111000001",
                      27 when "01111111000010",
                      27 when "01111111000011",
                      27 when "01111111000100",
                      27 when "01111111000101",
                      27 when "01111111000110",
                      27 when "01111111000111",
                      27 when "01111111001000",
                      27 when "01111111001001",
                      27 when "01111111001010",
                      27 when "01111111001011",
                      27 when "01111111001100",
                      27 when "01111111001101",
                      27 when "01111111001110",
                      27 when "01111111001111",
                      27 when "01111111010000",
                      27 when "01111111010001",
                      27 when "01111111010010",
                      27 when "01111111010011",
                      27 when "01111111010100",
                      27 when "01111111010101",
                      27 when "01111111010110",
                      27 when "01111111010111",
                      27 when "01111111011000",
                      27 when "01111111011001",
                      27 when "01111111011010",
                      27 when "01111111011011",
                      27 when "01111111011100",
                      27 when "01111111011101",
                      27 when "01111111011110",
                      27 when "01111111011111",
                      27 when "01111111100000",
                      27 when "01111111100001",
                      27 when "01111111100010",
                      27 when "01111111100011",
                      27 when "01111111100100",
                      27 when "01111111100101",
                      27 when "01111111100110",
                      27 when "01111111100111",
                      27 when "01111111101000",
                      27 when "01111111101001",
                      27 when "01111111101010",
                      27 when "01111111101011",
                      27 when "01111111101100",
                      27 when "01111111101101",
                      27 when "01111111101110",
                      27 when "01111111101111",
                      27 when "01111111110000",
                      27 when "01111111110001",
                      27 when "01111111110010",
                      27 when "01111111110011",
                      27 when "01111111110100",
                      27 when "01111111110101",
                      27 when "01111111110110",
                      27 when "01111111110111",
                      27 when "01111111111000",
                      27 when "01111111111001",
                      27 when "01111111111010",
                      27 when "01111111111011",
                      27 when "01111111111100",
                      27 when "01111111111101",
                      27 when "01111111111110",
                      27 when "01111111111111",
                      27 when "10000000000000",
                      27 when "10000000000001",
                      27 when "10000000000010",
                      27 when "10000000000011",
                      27 when "10000000000100",
                      27 when "10000000000101",
                      27 when "10000000000110",
                      27 when "10000000000111",
                      27 when "10000000001000",
                      27 when "10000000001001",
                      27 when "10000000001010",
                      27 when "10000000001011",
                      27 when "10000000001100",
                      27 when "10000000001101",
                      27 when "10000000001110",
                      27 when "10000000001111",
                      27 when "10000000010000",
                      27 when "10000000010001",
                      27 when "10000000010010",
                      27 when "10000000010011",
                      27 when "10000000010100",
                      27 when "10000000010101",
                      27 when "10000000010110",
                      27 when "10000000010111",
                      27 when "10000000011000",
                      27 when "10000000011001",
                      27 when "10000000011010",
                      27 when "10000000011011",
                      27 when "10000000011100",
                      27 when "10000000011101",
                      27 when "10000000011110",
                      27 when "10000000011111",
                      27 when "10000000100000",
                      27 when "10000000100001",
                      27 when "10000000100010",
                      27 when "10000000100011",
                      27 when "10000000100100",
                      27 when "10000000100101",
                      27 when "10000000100110",
                      27 when "10000000100111",
                      27 when "10000000101000",
                      27 when "10000000101001",
                      27 when "10000000101010",
                      27 when "10000000101011",
                      27 when "10000000101100",
                      27 when "10000000101101",
                      27 when "10000000101110",
                      27 when "10000000101111",
                      27 when "10000000110000",
                      27 when "10000000110001",
                      27 when "10000000110010",
                      27 when "10000000110011",
                      27 when "10000000110100",
                      27 when "10000000110101",
                      27 when "10000000110110",
                      27 when "10000000110111",
                      27 when "10000000111000",
                      27 when "10000000111001",
                      27 when "10000000111010",
                      27 when "10000000111011",
                      27 when "10000000111100",
                      27 when "10000000111101",
                      27 when "10000000111110",
                      27 when "10000000111111",
                      27 when "10000001000000",
                      27 when "10000001000001",
                      27 when "10000001000010",
                      27 when "10000001000011",
                      27 when "10000001000100",
                      27 when "10000001000101",
                      27 when "10000001000110",
                      27 when "10000001000111",
                      27 when "10000001001000",
                      27 when "10000001001001",
                      27 when "10000001001010",
                      27 when "10000001001011",
                      27 when "10000001001100",
                      27 when "10000001001101",
                      27 when "10000001001110",
                      27 when "10000001001111",
                      27 when "10000001010000",
                      27 when "10000001010001",
                      27 when "10000001010010",
                      27 when "10000001010011",
                      27 when "10000001010100",
                      27 when "10000001010101",
                      27 when "10000001010110",
                      27 when "10000001010111",
                      27 when "10000001011000",
                      27 when "10000001011001",
                      27 when "10000001011010",
                      27 when "10000001011011",
                      27 when "10000001011100",
                      27 when "10000001011101",
                      27 when "10000001011110",
                      27 when "10000001011111",
                      27 when "10000001100000",
                      27 when "10000001100001",
                      27 when "10000001100010",
                      27 when "10000001100011",
                      26 when "10000001100100",
                      26 when "10000001100101",
                      26 when "10000001100110",
                      26 when "10000001100111",
                      26 when "10000001101000",
                      26 when "10000001101001",
                      26 when "10000001101010",
                      26 when "10000001101011",
                      26 when "10000001101100",
                      26 when "10000001101101",
                      26 when "10000001101110",
                      26 when "10000001101111",
                      26 when "10000001110000",
                      26 when "10000001110001",
                      26 when "10000001110010",
                      26 when "10000001110011",
                      26 when "10000001110100",
                      26 when "10000001110101",
                      26 when "10000001110110",
                      26 when "10000001110111",
                      26 when "10000001111000",
                      26 when "10000001111001",
                      26 when "10000001111010",
                      26 when "10000001111011",
                      26 when "10000001111100",
                      26 when "10000001111101",
                      26 when "10000001111110",
                      26 when "10000001111111",
                      26 when "10000010000000",
                      26 when "10000010000001",
                      26 when "10000010000010",
                      26 when "10000010000011",
                      26 when "10000010000100",
                      26 when "10000010000101",
                      26 when "10000010000110",
                      26 when "10000010000111",
                      26 when "10000010001000",
                      26 when "10000010001001",
                      26 when "10000010001010",
                      26 when "10000010001011",
                      26 when "10000010001100",
                      26 when "10000010001101",
                      26 when "10000010001110",
                      26 when "10000010001111",
                      26 when "10000010010000",
                      26 when "10000010010001",
                      26 when "10000010010010",
                      26 when "10000010010011",
                      26 when "10000010010100",
                      26 when "10000010010101",
                      26 when "10000010010110",
                      26 when "10000010010111",
                      26 when "10000010011000",
                      26 when "10000010011001",
                      26 when "10000010011010",
                      26 when "10000010011011",
                      26 when "10000010011100",
                      26 when "10000010011101",
                      26 when "10000010011110",
                      26 when "10000010011111",
                      26 when "10000010100000",
                      26 when "10000010100001",
                      26 when "10000010100010",
                      26 when "10000010100011",
                      26 when "10000010100100",
                      26 when "10000010100101",
                      26 when "10000010100110",
                      26 when "10000010100111",
                      26 when "10000010101000",
                      26 when "10000010101001",
                      26 when "10000010101010",
                      26 when "10000010101011",
                      26 when "10000010101100",
                      26 when "10000010101101",
                      26 when "10000010101110",
                      26 when "10000010101111",
                      26 when "10000010110000",
                      26 when "10000010110001",
                      26 when "10000010110010",
                      26 when "10000010110011",
                      26 when "10000010110100",
                      26 when "10000010110101",
                      26 when "10000010110110",
                      26 when "10000010110111",
                      26 when "10000010111000",
                      26 when "10000010111001",
                      26 when "10000010111010",
                      26 when "10000010111011",
                      26 when "10000010111100",
                      26 when "10000010111101",
                      26 when "10000010111110",
                      26 when "10000010111111",
                      26 when "10000011000000",
                      26 when "10000011000001",
                      26 when "10000011000010",
                      26 when "10000011000011",
                      26 when "10000011000100",
                      26 when "10000011000101",
                      26 when "10000011000110",
                      26 when "10000011000111",
                      26 when "10000011001000",
                      26 when "10000011001001",
                      26 when "10000011001010",
                      26 when "10000011001011",
                      26 when "10000011001100",
                      26 when "10000011001101",
                      26 when "10000011001110",
                      26 when "10000011001111",
                      26 when "10000011010000",
                      26 when "10000011010001",
                      26 when "10000011010010",
                      26 when "10000011010011",
                      26 when "10000011010100",
                      26 when "10000011010101",
                      26 when "10000011010110",
                      26 when "10000011010111",
                      26 when "10000011011000",
                      26 when "10000011011001",
                      26 when "10000011011010",
                      26 when "10000011011011",
                      26 when "10000011011100",
                      26 when "10000011011101",
                      26 when "10000011011110",
                      26 when "10000011011111",
                      26 when "10000011100000",
                      26 when "10000011100001",
                      26 when "10000011100010",
                      26 when "10000011100011",
                      26 when "10000011100100",
                      26 when "10000011100101",
                      26 when "10000011100110",
                      26 when "10000011100111",
                      26 when "10000011101000",
                      26 when "10000011101001",
                      26 when "10000011101010",
                      26 when "10000011101011",
                      26 when "10000011101100",
                      26 when "10000011101101",
                      26 when "10000011101110",
                      26 when "10000011101111",
                      26 when "10000011110000",
                      26 when "10000011110001",
                      26 when "10000011110010",
                      26 when "10000011110011",
                      26 when "10000011110100",
                      26 when "10000011110101",
                      26 when "10000011110110",
                      26 when "10000011110111",
                      26 when "10000011111000",
                      26 when "10000011111001",
                      26 when "10000011111010",
                      26 when "10000011111011",
                      26 when "10000011111100",
                      26 when "10000011111101",
                      26 when "10000011111110",
                      26 when "10000011111111",
                      26 when "10000100000000",
                      26 when "10000100000001",
                      26 when "10000100000010",
                      26 when "10000100000011",
                      26 when "10000100000100",
                      26 when "10000100000101",
                      26 when "10000100000110",
                      26 when "10000100000111",
                      26 when "10000100001000",
                      26 when "10000100001001",
                      26 when "10000100001010",
                      26 when "10000100001011",
                      26 when "10000100001100",
                      26 when "10000100001101",
                      26 when "10000100001110",
                      26 when "10000100001111",
                      26 when "10000100010000",
                      26 when "10000100010001",
                      26 when "10000100010010",
                      26 when "10000100010011",
                      26 when "10000100010100",
                      26 when "10000100010101",
                      26 when "10000100010110",
                      26 when "10000100010111",
                      26 when "10000100011000",
                      26 when "10000100011001",
                      26 when "10000100011010",
                      26 when "10000100011011",
                      26 when "10000100011100",
                      26 when "10000100011101",
                      26 when "10000100011110",
                      26 when "10000100011111",
                      26 when "10000100100000",
                      26 when "10000100100001",
                      26 when "10000100100010",
                      26 when "10000100100011",
                      26 when "10000100100100",
                      26 when "10000100100101",
                      26 when "10000100100110",
                      26 when "10000100100111",
                      26 when "10000100101000",
                      26 when "10000100101001",
                      26 when "10000100101010",
                      26 when "10000100101011",
                      26 when "10000100101100",
                      26 when "10000100101101",
                      26 when "10000100101110",
                      26 when "10000100101111",
                      26 when "10000100110000",
                      26 when "10000100110001",
                      26 when "10000100110010",
                      26 when "10000100110011",
                      26 when "10000100110100",
                      26 when "10000100110101",
                      26 when "10000100110110",
                      26 when "10000100110111",
                      26 when "10000100111000",
                      26 when "10000100111001",
                      26 when "10000100111010",
                      26 when "10000100111011",
                      26 when "10000100111100",
                      26 when "10000100111101",
                      26 when "10000100111110",
                      26 when "10000100111111",
                      26 when "10000101000000",
                      26 when "10000101000001",
                      26 when "10000101000010",
                      26 when "10000101000011",
                      26 when "10000101000100",
                      26 when "10000101000101",
                      26 when "10000101000110",
                      26 when "10000101000111",
                      26 when "10000101001000",
                      26 when "10000101001001",
                      26 when "10000101001010",
                      26 when "10000101001011",
                      26 when "10000101001100",
                      26 when "10000101001101",
                      26 when "10000101001110",
                      26 when "10000101001111",
                      26 when "10000101010000",
                      26 when "10000101010001",
                      26 when "10000101010010",
                      26 when "10000101010011",
                      26 when "10000101010100",
                      26 when "10000101010101",
                      26 when "10000101010110",
                      26 when "10000101010111",
                      26 when "10000101011000",
                      26 when "10000101011001",
                      26 when "10000101011010",
                      26 when "10000101011011",
                      26 when "10000101011100",
                      26 when "10000101011101",
                      26 when "10000101011110",
                      26 when "10000101011111",
                      26 when "10000101100000",
                      26 when "10000101100001",
                      26 when "10000101100010",
                      26 when "10000101100011",
                      26 when "10000101100100",
                      26 when "10000101100101",
                      26 when "10000101100110",
                      26 when "10000101100111",
                      26 when "10000101101000",
                      26 when "10000101101001",
                      26 when "10000101101010",
                      26 when "10000101101011",
                      26 when "10000101101100",
                      26 when "10000101101101",
                      26 when "10000101101110",
                      26 when "10000101101111",
                      26 when "10000101110000",
                      26 when "10000101110001",
                      26 when "10000101110010",
                      26 when "10000101110011",
                      26 when "10000101110100",
                      26 when "10000101110101",
                      26 when "10000101110110",
                      26 when "10000101110111",
                      26 when "10000101111000",
                      26 when "10000101111001",
                      26 when "10000101111010",
                      26 when "10000101111011",
                      26 when "10000101111100",
                      26 when "10000101111101",
                      26 when "10000101111110",
                      26 when "10000101111111",
                      26 when "10000110000000",
                      26 when "10000110000001",
                      26 when "10000110000010",
                      26 when "10000110000011",
                      26 when "10000110000100",
                      26 when "10000110000101",
                      26 when "10000110000110",
                      26 when "10000110000111",
                      26 when "10000110001000",
                      26 when "10000110001001",
                      26 when "10000110001010",
                      26 when "10000110001011",
                      26 when "10000110001100",
                      26 when "10000110001101",
                      26 when "10000110001110",
                      26 when "10000110001111",
                      26 when "10000110010000",
                      26 when "10000110010001",
                      26 when "10000110010010",
                      26 when "10000110010011",
                      26 when "10000110010100",
                      26 when "10000110010101",
                      26 when "10000110010110",
                      26 when "10000110010111",
                      26 when "10000110011000",
                      26 when "10000110011001",
                      26 when "10000110011010",
                      26 when "10000110011011",
                      26 when "10000110011100",
                      26 when "10000110011101",
                      26 when "10000110011110",
                      26 when "10000110011111",
                      26 when "10000110100000",
                      26 when "10000110100001",
                      26 when "10000110100010",
                      26 when "10000110100011",
                      26 when "10000110100100",
                      26 when "10000110100101",
                      26 when "10000110100110",
                      26 when "10000110100111",
                      26 when "10000110101000",
                      25 when "10000110101001",
                      25 when "10000110101010",
                      25 when "10000110101011",
                      25 when "10000110101100",
                      25 when "10000110101101",
                      25 when "10000110101110",
                      25 when "10000110101111",
                      25 when "10000110110000",
                      25 when "10000110110001",
                      25 when "10000110110010",
                      25 when "10000110110011",
                      25 when "10000110110100",
                      25 when "10000110110101",
                      25 when "10000110110110",
                      25 when "10000110110111",
                      25 when "10000110111000",
                      25 when "10000110111001",
                      25 when "10000110111010",
                      25 when "10000110111011",
                      25 when "10000110111100",
                      25 when "10000110111101",
                      25 when "10000110111110",
                      25 when "10000110111111",
                      25 when "10000111000000",
                      25 when "10000111000001",
                      25 when "10000111000010",
                      25 when "10000111000011",
                      25 when "10000111000100",
                      25 when "10000111000101",
                      25 when "10000111000110",
                      25 when "10000111000111",
                      25 when "10000111001000",
                      25 when "10000111001001",
                      25 when "10000111001010",
                      25 when "10000111001011",
                      25 when "10000111001100",
                      25 when "10000111001101",
                      25 when "10000111001110",
                      25 when "10000111001111",
                      25 when "10000111010000",
                      25 when "10000111010001",
                      25 when "10000111010010",
                      25 when "10000111010011",
                      25 when "10000111010100",
                      25 when "10000111010101",
                      25 when "10000111010110",
                      25 when "10000111010111",
                      25 when "10000111011000",
                      25 when "10000111011001",
                      25 when "10000111011010",
                      25 when "10000111011011",
                      25 when "10000111011100",
                      25 when "10000111011101",
                      25 when "10000111011110",
                      25 when "10000111011111",
                      25 when "10000111100000",
                      25 when "10000111100001",
                      25 when "10000111100010",
                      25 when "10000111100011",
                      25 when "10000111100100",
                      25 when "10000111100101",
                      25 when "10000111100110",
                      25 when "10000111100111",
                      25 when "10000111101000",
                      25 when "10000111101001",
                      25 when "10000111101010",
                      25 when "10000111101011",
                      25 when "10000111101100",
                      25 when "10000111101101",
                      25 when "10000111101110",
                      25 when "10000111101111",
                      25 when "10000111110000",
                      25 when "10000111110001",
                      25 when "10000111110010",
                      25 when "10000111110011",
                      25 when "10000111110100",
                      25 when "10000111110101",
                      25 when "10000111110110",
                      25 when "10000111110111",
                      25 when "10000111111000",
                      25 when "10000111111001",
                      25 when "10000111111010",
                      25 when "10000111111011",
                      25 when "10000111111100",
                      25 when "10000111111101",
                      25 when "10000111111110",
                      25 when "10000111111111",
                      25 when "10001000000000",
                      25 when "10001000000001",
                      25 when "10001000000010",
                      25 when "10001000000011",
                      25 when "10001000000100",
                      25 when "10001000000101",
                      25 when "10001000000110",
                      25 when "10001000000111",
                      25 when "10001000001000",
                      25 when "10001000001001",
                      25 when "10001000001010",
                      25 when "10001000001011",
                      25 when "10001000001100",
                      25 when "10001000001101",
                      25 when "10001000001110",
                      25 when "10001000001111",
                      25 when "10001000010000",
                      25 when "10001000010001",
                      25 when "10001000010010",
                      25 when "10001000010011",
                      25 when "10001000010100",
                      25 when "10001000010101",
                      25 when "10001000010110",
                      25 when "10001000010111",
                      25 when "10001000011000",
                      25 when "10001000011001",
                      25 when "10001000011010",
                      25 when "10001000011011",
                      25 when "10001000011100",
                      25 when "10001000011101",
                      25 when "10001000011110",
                      25 when "10001000011111",
                      25 when "10001000100000",
                      25 when "10001000100001",
                      25 when "10001000100010",
                      25 when "10001000100011",
                      25 when "10001000100100",
                      25 when "10001000100101",
                      25 when "10001000100110",
                      25 when "10001000100111",
                      25 when "10001000101000",
                      25 when "10001000101001",
                      25 when "10001000101010",
                      25 when "10001000101011",
                      25 when "10001000101100",
                      25 when "10001000101101",
                      25 when "10001000101110",
                      25 when "10001000101111",
                      25 when "10001000110000",
                      25 when "10001000110001",
                      25 when "10001000110010",
                      25 when "10001000110011",
                      25 when "10001000110100",
                      25 when "10001000110101",
                      25 when "10001000110110",
                      25 when "10001000110111",
                      25 when "10001000111000",
                      25 when "10001000111001",
                      25 when "10001000111010",
                      25 when "10001000111011",
                      25 when "10001000111100",
                      25 when "10001000111101",
                      25 when "10001000111110",
                      25 when "10001000111111",
                      25 when "10001001000000",
                      25 when "10001001000001",
                      25 when "10001001000010",
                      25 when "10001001000011",
                      25 when "10001001000100",
                      25 when "10001001000101",
                      25 when "10001001000110",
                      25 when "10001001000111",
                      25 when "10001001001000",
                      25 when "10001001001001",
                      25 when "10001001001010",
                      25 when "10001001001011",
                      25 when "10001001001100",
                      25 when "10001001001101",
                      25 when "10001001001110",
                      25 when "10001001001111",
                      25 when "10001001010000",
                      25 when "10001001010001",
                      25 when "10001001010010",
                      25 when "10001001010011",
                      25 when "10001001010100",
                      25 when "10001001010101",
                      25 when "10001001010110",
                      25 when "10001001010111",
                      25 when "10001001011000",
                      25 when "10001001011001",
                      25 when "10001001011010",
                      25 when "10001001011011",
                      25 when "10001001011100",
                      25 when "10001001011101",
                      25 when "10001001011110",
                      25 when "10001001011111",
                      25 when "10001001100000",
                      25 when "10001001100001",
                      25 when "10001001100010",
                      25 when "10001001100011",
                      25 when "10001001100100",
                      25 when "10001001100101",
                      25 when "10001001100110",
                      25 when "10001001100111",
                      25 when "10001001101000",
                      25 when "10001001101001",
                      25 when "10001001101010",
                      25 when "10001001101011",
                      25 when "10001001101100",
                      25 when "10001001101101",
                      25 when "10001001101110",
                      25 when "10001001101111",
                      25 when "10001001110000",
                      25 when "10001001110001",
                      25 when "10001001110010",
                      25 when "10001001110011",
                      25 when "10001001110100",
                      25 when "10001001110101",
                      25 when "10001001110110",
                      25 when "10001001110111",
                      25 when "10001001111000",
                      25 when "10001001111001",
                      25 when "10001001111010",
                      25 when "10001001111011",
                      25 when "10001001111100",
                      25 when "10001001111101",
                      25 when "10001001111110",
                      25 when "10001001111111",
                      25 when "10001010000000",
                      25 when "10001010000001",
                      25 when "10001010000010",
                      25 when "10001010000011",
                      25 when "10001010000100",
                      25 when "10001010000101",
                      25 when "10001010000110",
                      25 when "10001010000111",
                      25 when "10001010001000",
                      25 when "10001010001001",
                      25 when "10001010001010",
                      25 when "10001010001011",
                      25 when "10001010001100",
                      25 when "10001010001101",
                      25 when "10001010001110",
                      25 when "10001010001111",
                      25 when "10001010010000",
                      25 when "10001010010001",
                      25 when "10001010010010",
                      25 when "10001010010011",
                      25 when "10001010010100",
                      25 when "10001010010101",
                      25 when "10001010010110",
                      25 when "10001010010111",
                      25 when "10001010011000",
                      25 when "10001010011001",
                      25 when "10001010011010",
                      25 when "10001010011011",
                      25 when "10001010011100",
                      25 when "10001010011101",
                      25 when "10001010011110",
                      25 when "10001010011111",
                      25 when "10001010100000",
                      25 when "10001010100001",
                      25 when "10001010100010",
                      25 when "10001010100011",
                      25 when "10001010100100",
                      25 when "10001010100101",
                      25 when "10001010100110",
                      25 when "10001010100111",
                      25 when "10001010101000",
                      25 when "10001010101001",
                      25 when "10001010101010",
                      25 when "10001010101011",
                      25 when "10001010101100",
                      25 when "10001010101101",
                      25 when "10001010101110",
                      25 when "10001010101111",
                      25 when "10001010110000",
                      25 when "10001010110001",
                      25 when "10001010110010",
                      25 when "10001010110011",
                      25 when "10001010110100",
                      25 when "10001010110101",
                      25 when "10001010110110",
                      25 when "10001010110111",
                      25 when "10001010111000",
                      25 when "10001010111001",
                      25 when "10001010111010",
                      25 when "10001010111011",
                      25 when "10001010111100",
                      25 when "10001010111101",
                      25 when "10001010111110",
                      25 when "10001010111111",
                      25 when "10001011000000",
                      25 when "10001011000001",
                      25 when "10001011000010",
                      25 when "10001011000011",
                      25 when "10001011000100",
                      25 when "10001011000101",
                      25 when "10001011000110",
                      25 when "10001011000111",
                      25 when "10001011001000",
                      25 when "10001011001001",
                      25 when "10001011001010",
                      25 when "10001011001011",
                      25 when "10001011001100",
                      25 when "10001011001101",
                      25 when "10001011001110",
                      25 when "10001011001111",
                      25 when "10001011010000",
                      25 when "10001011010001",
                      25 when "10001011010010",
                      25 when "10001011010011",
                      25 when "10001011010100",
                      25 when "10001011010101",
                      25 when "10001011010110",
                      25 when "10001011010111",
                      25 when "10001011011000",
                      25 when "10001011011001",
                      25 when "10001011011010",
                      25 when "10001011011011",
                      25 when "10001011011100",
                      25 when "10001011011101",
                      25 when "10001011011110",
                      25 when "10001011011111",
                      25 when "10001011100000",
                      25 when "10001011100001",
                      25 when "10001011100010",
                      25 when "10001011100011",
                      25 when "10001011100100",
                      25 when "10001011100101",
                      25 when "10001011100110",
                      25 when "10001011100111",
                      25 when "10001011101000",
                      25 when "10001011101001",
                      25 when "10001011101010",
                      25 when "10001011101011",
                      25 when "10001011101100",
                      25 when "10001011101101",
                      25 when "10001011101110",
                      25 when "10001011101111",
                      25 when "10001011110000",
                      25 when "10001011110001",
                      25 when "10001011110010",
                      25 when "10001011110011",
                      25 when "10001011110100",
                      25 when "10001011110101",
                      25 when "10001011110110",
                      25 when "10001011110111",
                      25 when "10001011111000",
                      25 when "10001011111001",
                      25 when "10001011111010",
                      25 when "10001011111011",
                      25 when "10001011111100",
                      25 when "10001011111101",
                      25 when "10001011111110",
                      25 when "10001011111111",
                      25 when "10001100000000",
                      25 when "10001100000001",
                      25 when "10001100000010",
                      25 when "10001100000011",
                      25 when "10001100000100",
                      25 when "10001100000101",
                      25 when "10001100000110",
                      25 when "10001100000111",
                      25 when "10001100001000",
                      24 when "10001100001001",
                      24 when "10001100001010",
                      24 when "10001100001011",
                      24 when "10001100001100",
                      24 when "10001100001101",
                      24 when "10001100001110",
                      24 when "10001100001111",
                      24 when "10001100010000",
                      24 when "10001100010001",
                      24 when "10001100010010",
                      24 when "10001100010011",
                      24 when "10001100010100",
                      24 when "10001100010101",
                      24 when "10001100010110",
                      24 when "10001100010111",
                      24 when "10001100011000",
                      24 when "10001100011001",
                      24 when "10001100011010",
                      24 when "10001100011011",
                      24 when "10001100011100",
                      24 when "10001100011101",
                      24 when "10001100011110",
                      24 when "10001100011111",
                      24 when "10001100100000",
                      24 when "10001100100001",
                      24 when "10001100100010",
                      24 when "10001100100011",
                      24 when "10001100100100",
                      24 when "10001100100101",
                      24 when "10001100100110",
                      24 when "10001100100111",
                      24 when "10001100101000",
                      24 when "10001100101001",
                      24 when "10001100101010",
                      24 when "10001100101011",
                      24 when "10001100101100",
                      24 when "10001100101101",
                      24 when "10001100101110",
                      24 when "10001100101111",
                      24 when "10001100110000",
                      24 when "10001100110001",
                      24 when "10001100110010",
                      24 when "10001100110011",
                      24 when "10001100110100",
                      24 when "10001100110101",
                      24 when "10001100110110",
                      24 when "10001100110111",
                      24 when "10001100111000",
                      24 when "10001100111001",
                      24 when "10001100111010",
                      24 when "10001100111011",
                      24 when "10001100111100",
                      24 when "10001100111101",
                      24 when "10001100111110",
                      24 when "10001100111111",
                      24 when "10001101000000",
                      24 when "10001101000001",
                      24 when "10001101000010",
                      24 when "10001101000011",
                      24 when "10001101000100",
                      24 when "10001101000101",
                      24 when "10001101000110",
                      24 when "10001101000111",
                      24 when "10001101001000",
                      24 when "10001101001001",
                      24 when "10001101001010",
                      24 when "10001101001011",
                      24 when "10001101001100",
                      24 when "10001101001101",
                      24 when "10001101001110",
                      24 when "10001101001111",
                      24 when "10001101010000",
                      24 when "10001101010001",
                      24 when "10001101010010",
                      24 when "10001101010011",
                      24 when "10001101010100",
                      24 when "10001101010101",
                      24 when "10001101010110",
                      24 when "10001101010111",
                      24 when "10001101011000",
                      24 when "10001101011001",
                      24 when "10001101011010",
                      24 when "10001101011011",
                      24 when "10001101011100",
                      24 when "10001101011101",
                      24 when "10001101011110",
                      24 when "10001101011111",
                      24 when "10001101100000",
                      24 when "10001101100001",
                      24 when "10001101100010",
                      24 when "10001101100011",
                      24 when "10001101100100",
                      24 when "10001101100101",
                      24 when "10001101100110",
                      24 when "10001101100111",
                      24 when "10001101101000",
                      24 when "10001101101001",
                      24 when "10001101101010",
                      24 when "10001101101011",
                      24 when "10001101101100",
                      24 when "10001101101101",
                      24 when "10001101101110",
                      24 when "10001101101111",
                      24 when "10001101110000",
                      24 when "10001101110001",
                      24 when "10001101110010",
                      24 when "10001101110011",
                      24 when "10001101110100",
                      24 when "10001101110101",
                      24 when "10001101110110",
                      24 when "10001101110111",
                      24 when "10001101111000",
                      24 when "10001101111001",
                      24 when "10001101111010",
                      24 when "10001101111011",
                      24 when "10001101111100",
                      24 when "10001101111101",
                      24 when "10001101111110",
                      24 when "10001101111111",
                      24 when "10001110000000",
                      24 when "10001110000001",
                      24 when "10001110000010",
                      24 when "10001110000011",
                      24 when "10001110000100",
                      24 when "10001110000101",
                      24 when "10001110000110",
                      24 when "10001110000111",
                      24 when "10001110001000",
                      24 when "10001110001001",
                      24 when "10001110001010",
                      24 when "10001110001011",
                      24 when "10001110001100",
                      24 when "10001110001101",
                      24 when "10001110001110",
                      24 when "10001110001111",
                      24 when "10001110010000",
                      24 when "10001110010001",
                      24 when "10001110010010",
                      24 when "10001110010011",
                      24 when "10001110010100",
                      24 when "10001110010101",
                      24 when "10001110010110",
                      24 when "10001110010111",
                      24 when "10001110011000",
                      24 when "10001110011001",
                      24 when "10001110011010",
                      24 when "10001110011011",
                      24 when "10001110011100",
                      24 when "10001110011101",
                      24 when "10001110011110",
                      24 when "10001110011111",
                      24 when "10001110100000",
                      24 when "10001110100001",
                      24 when "10001110100010",
                      24 when "10001110100011",
                      24 when "10001110100100",
                      24 when "10001110100101",
                      24 when "10001110100110",
                      24 when "10001110100111",
                      24 when "10001110101000",
                      24 when "10001110101001",
                      24 when "10001110101010",
                      24 when "10001110101011",
                      24 when "10001110101100",
                      24 when "10001110101101",
                      24 when "10001110101110",
                      24 when "10001110101111",
                      24 when "10001110110000",
                      24 when "10001110110001",
                      24 when "10001110110010",
                      24 when "10001110110011",
                      24 when "10001110110100",
                      24 when "10001110110101",
                      24 when "10001110110110",
                      24 when "10001110110111",
                      24 when "10001110111000",
                      24 when "10001110111001",
                      24 when "10001110111010",
                      24 when "10001110111011",
                      24 when "10001110111100",
                      24 when "10001110111101",
                      24 when "10001110111110",
                      24 when "10001110111111",
                      24 when "10001111000000",
                      24 when "10001111000001",
                      24 when "10001111000010",
                      24 when "10001111000011",
                      24 when "10001111000100",
                      24 when "10001111000101",
                      24 when "10001111000110",
                      24 when "10001111000111",
                      24 when "10001111001000",
                      24 when "10001111001001",
                      24 when "10001111001010",
                      24 when "10001111001011",
                      24 when "10001111001100",
                      24 when "10001111001101",
                      24 when "10001111001110",
                      24 when "10001111001111",
                      24 when "10001111010000",
                      24 when "10001111010001",
                      24 when "10001111010010",
                      24 when "10001111010011",
                      24 when "10001111010100",
                      24 when "10001111010101",
                      24 when "10001111010110",
                      24 when "10001111010111",
                      24 when "10001111011000",
                      24 when "10001111011001",
                      24 when "10001111011010",
                      24 when "10001111011011",
                      24 when "10001111011100",
                      24 when "10001111011101",
                      24 when "10001111011110",
                      24 when "10001111011111",
                      24 when "10001111100000",
                      24 when "10001111100001",
                      24 when "10001111100010",
                      24 when "10001111100011",
                      24 when "10001111100100",
                      24 when "10001111100101",
                      24 when "10001111100110",
                      24 when "10001111100111",
                      24 when "10001111101000",
                      24 when "10001111101001",
                      24 when "10001111101010",
                      24 when "10001111101011",
                      24 when "10001111101100",
                      24 when "10001111101101",
                      24 when "10001111101110",
                      24 when "10001111101111",
                      24 when "10001111110000",
                      24 when "10001111110001",
                      24 when "10001111110010",
                      24 when "10001111110011",
                      24 when "10001111110100",
                      24 when "10001111110101",
                      24 when "10001111110110",
                      24 when "10001111110111",
                      24 when "10001111111000",
                      24 when "10001111111001",
                      24 when "10001111111010",
                      24 when "10001111111011",
                      24 when "10001111111100",
                      24 when "10001111111101",
                      24 when "10001111111110",
                      24 when "10001111111111",
                      24 when "10010000000000",
                      24 when "10010000000001",
                      24 when "10010000000010",
                      24 when "10010000000011",
                      24 when "10010000000100",
                      24 when "10010000000101",
                      24 when "10010000000110",
                      24 when "10010000000111",
                      24 when "10010000001000",
                      24 when "10010000001001",
                      24 when "10010000001010",
                      24 when "10010000001011",
                      24 when "10010000001100",
                      24 when "10010000001101",
                      24 when "10010000001110",
                      24 when "10010000001111",
                      24 when "10010000010000",
                      24 when "10010000010001",
                      24 when "10010000010010",
                      24 when "10010000010011",
                      24 when "10010000010100",
                      24 when "10010000010101",
                      24 when "10010000010110",
                      24 when "10010000010111",
                      24 when "10010000011000",
                      24 when "10010000011001",
                      24 when "10010000011010",
                      24 when "10010000011011",
                      24 when "10010000011100",
                      24 when "10010000011101",
                      24 when "10010000011110",
                      24 when "10010000011111",
                      24 when "10010000100000",
                      24 when "10010000100001",
                      24 when "10010000100010",
                      24 when "10010000100011",
                      24 when "10010000100100",
                      24 when "10010000100101",
                      24 when "10010000100110",
                      24 when "10010000100111",
                      24 when "10010000101000",
                      24 when "10010000101001",
                      24 when "10010000101010",
                      24 when "10010000101011",
                      24 when "10010000101100",
                      24 when "10010000101101",
                      24 when "10010000101110",
                      24 when "10010000101111",
                      24 when "10010000110000",
                      24 when "10010000110001",
                      24 when "10010000110010",
                      24 when "10010000110011",
                      24 when "10010000110100",
                      24 when "10010000110101",
                      24 when "10010000110110",
                      24 when "10010000110111",
                      24 when "10010000111000",
                      24 when "10010000111001",
                      24 when "10010000111010",
                      24 when "10010000111011",
                      24 when "10010000111100",
                      24 when "10010000111101",
                      24 when "10010000111110",
                      24 when "10010000111111",
                      24 when "10010001000000",
                      24 when "10010001000001",
                      24 when "10010001000010",
                      24 when "10010001000011",
                      24 when "10010001000100",
                      24 when "10010001000101",
                      24 when "10010001000110",
                      24 when "10010001000111",
                      24 when "10010001001000",
                      24 when "10010001001001",
                      24 when "10010001001010",
                      24 when "10010001001011",
                      24 when "10010001001100",
                      24 when "10010001001101",
                      24 when "10010001001110",
                      24 when "10010001001111",
                      24 when "10010001010000",
                      24 when "10010001010001",
                      24 when "10010001010010",
                      24 when "10010001010011",
                      24 when "10010001010100",
                      24 when "10010001010101",
                      24 when "10010001010110",
                      24 when "10010001010111",
                      24 when "10010001011000",
                      24 when "10010001011001",
                      24 when "10010001011010",
                      24 when "10010001011011",
                      24 when "10010001011100",
                      24 when "10010001011101",
                      24 when "10010001011110",
                      24 when "10010001011111",
                      24 when "10010001100000",
                      24 when "10010001100001",
                      24 when "10010001100010",
                      24 when "10010001100011",
                      24 when "10010001100100",
                      24 when "10010001100101",
                      24 when "10010001100110",
                      24 when "10010001100111",
                      24 when "10010001101000",
                      24 when "10010001101001",
                      24 when "10010001101010",
                      24 when "10010001101011",
                      24 when "10010001101100",
                      24 when "10010001101101",
                      24 when "10010001101110",
                      24 when "10010001101111",
                      24 when "10010001110000",
                      24 when "10010001110001",
                      24 when "10010001110010",
                      24 when "10010001110011",
                      24 when "10010001110100",
                      24 when "10010001110101",
                      24 when "10010001110110",
                      24 when "10010001110111",
                      24 when "10010001111000",
                      24 when "10010001111001",
                      24 when "10010001111010",
                      24 when "10010001111011",
                      24 when "10010001111100",
                      24 when "10010001111101",
                      24 when "10010001111110",
                      24 when "10010001111111",
                      24 when "10010010000000",
                      24 when "10010010000001",
                      24 when "10010010000010",
                      24 when "10010010000011",
                      24 when "10010010000100",
                      24 when "10010010000101",
                      24 when "10010010000110",
                      23 when "10010010000111",
                      23 when "10010010001000",
                      23 when "10010010001001",
                      23 when "10010010001010",
                      23 when "10010010001011",
                      23 when "10010010001100",
                      23 when "10010010001101",
                      23 when "10010010001110",
                      23 when "10010010001111",
                      23 when "10010010010000",
                      23 when "10010010010001",
                      23 when "10010010010010",
                      23 when "10010010010011",
                      23 when "10010010010100",
                      23 when "10010010010101",
                      23 when "10010010010110",
                      23 when "10010010010111",
                      23 when "10010010011000",
                      23 when "10010010011001",
                      23 when "10010010011010",
                      23 when "10010010011011",
                      23 when "10010010011100",
                      23 when "10010010011101",
                      23 when "10010010011110",
                      23 when "10010010011111",
                      23 when "10010010100000",
                      23 when "10010010100001",
                      23 when "10010010100010",
                      23 when "10010010100011",
                      23 when "10010010100100",
                      23 when "10010010100101",
                      23 when "10010010100110",
                      23 when "10010010100111",
                      23 when "10010010101000",
                      23 when "10010010101001",
                      23 when "10010010101010",
                      23 when "10010010101011",
                      23 when "10010010101100",
                      23 when "10010010101101",
                      23 when "10010010101110",
                      23 when "10010010101111",
                      23 when "10010010110000",
                      23 when "10010010110001",
                      23 when "10010010110010",
                      23 when "10010010110011",
                      23 when "10010010110100",
                      23 when "10010010110101",
                      23 when "10010010110110",
                      23 when "10010010110111",
                      23 when "10010010111000",
                      23 when "10010010111001",
                      23 when "10010010111010",
                      23 when "10010010111011",
                      23 when "10010010111100",
                      23 when "10010010111101",
                      23 when "10010010111110",
                      23 when "10010010111111",
                      23 when "10010011000000",
                      23 when "10010011000001",
                      23 when "10010011000010",
                      23 when "10010011000011",
                      23 when "10010011000100",
                      23 when "10010011000101",
                      23 when "10010011000110",
                      23 when "10010011000111",
                      23 when "10010011001000",
                      23 when "10010011001001",
                      23 when "10010011001010",
                      23 when "10010011001011",
                      23 when "10010011001100",
                      23 when "10010011001101",
                      23 when "10010011001110",
                      23 when "10010011001111",
                      23 when "10010011010000",
                      23 when "10010011010001",
                      23 when "10010011010010",
                      23 when "10010011010011",
                      23 when "10010011010100",
                      23 when "10010011010101",
                      23 when "10010011010110",
                      23 when "10010011010111",
                      23 when "10010011011000",
                      23 when "10010011011001",
                      23 when "10010011011010",
                      23 when "10010011011011",
                      23 when "10010011011100",
                      23 when "10010011011101",
                      23 when "10010011011110",
                      23 when "10010011011111",
                      23 when "10010011100000",
                      23 when "10010011100001",
                      23 when "10010011100010",
                      23 when "10010011100011",
                      23 when "10010011100100",
                      23 when "10010011100101",
                      23 when "10010011100110",
                      23 when "10010011100111",
                      23 when "10010011101000",
                      23 when "10010011101001",
                      23 when "10010011101010",
                      23 when "10010011101011",
                      23 when "10010011101100",
                      23 when "10010011101101",
                      23 when "10010011101110",
                      23 when "10010011101111",
                      23 when "10010011110000",
                      23 when "10010011110001",
                      23 when "10010011110010",
                      23 when "10010011110011",
                      23 when "10010011110100",
                      23 when "10010011110101",
                      23 when "10010011110110",
                      23 when "10010011110111",
                      23 when "10010011111000",
                      23 when "10010011111001",
                      23 when "10010011111010",
                      23 when "10010011111011",
                      23 when "10010011111100",
                      23 when "10010011111101",
                      23 when "10010011111110",
                      23 when "10010011111111",
                      23 when "10010100000000",
                      23 when "10010100000001",
                      23 when "10010100000010",
                      23 when "10010100000011",
                      23 when "10010100000100",
                      23 when "10010100000101",
                      23 when "10010100000110",
                      23 when "10010100000111",
                      23 when "10010100001000",
                      23 when "10010100001001",
                      23 when "10010100001010",
                      23 when "10010100001011",
                      23 when "10010100001100",
                      23 when "10010100001101",
                      23 when "10010100001110",
                      23 when "10010100001111",
                      23 when "10010100010000",
                      23 when "10010100010001",
                      23 when "10010100010010",
                      23 when "10010100010011",
                      23 when "10010100010100",
                      23 when "10010100010101",
                      23 when "10010100010110",
                      23 when "10010100010111",
                      23 when "10010100011000",
                      23 when "10010100011001",
                      23 when "10010100011010",
                      23 when "10010100011011",
                      23 when "10010100011100",
                      23 when "10010100011101",
                      23 when "10010100011110",
                      23 when "10010100011111",
                      23 when "10010100100000",
                      23 when "10010100100001",
                      23 when "10010100100010",
                      23 when "10010100100011",
                      23 when "10010100100100",
                      23 when "10010100100101",
                      23 when "10010100100110",
                      23 when "10010100100111",
                      23 when "10010100101000",
                      23 when "10010100101001",
                      23 when "10010100101010",
                      23 when "10010100101011",
                      23 when "10010100101100",
                      23 when "10010100101101",
                      23 when "10010100101110",
                      23 when "10010100101111",
                      23 when "10010100110000",
                      23 when "10010100110001",
                      23 when "10010100110010",
                      23 when "10010100110011",
                      23 when "10010100110100",
                      23 when "10010100110101",
                      23 when "10010100110110",
                      23 when "10010100110111",
                      23 when "10010100111000",
                      23 when "10010100111001",
                      23 when "10010100111010",
                      23 when "10010100111011",
                      23 when "10010100111100",
                      23 when "10010100111101",
                      23 when "10010100111110",
                      23 when "10010100111111",
                      23 when "10010101000000",
                      23 when "10010101000001",
                      23 when "10010101000010",
                      23 when "10010101000011",
                      23 when "10010101000100",
                      23 when "10010101000101",
                      23 when "10010101000110",
                      23 when "10010101000111",
                      23 when "10010101001000",
                      23 when "10010101001001",
                      23 when "10010101001010",
                      23 when "10010101001011",
                      23 when "10010101001100",
                      23 when "10010101001101",
                      23 when "10010101001110",
                      23 when "10010101001111",
                      23 when "10010101010000",
                      23 when "10010101010001",
                      23 when "10010101010010",
                      23 when "10010101010011",
                      23 when "10010101010100",
                      23 when "10010101010101",
                      23 when "10010101010110",
                      23 when "10010101010111",
                      23 when "10010101011000",
                      23 when "10010101011001",
                      23 when "10010101011010",
                      23 when "10010101011011",
                      23 when "10010101011100",
                      23 when "10010101011101",
                      23 when "10010101011110",
                      23 when "10010101011111",
                      23 when "10010101100000",
                      23 when "10010101100001",
                      23 when "10010101100010",
                      23 when "10010101100011",
                      23 when "10010101100100",
                      23 when "10010101100101",
                      23 when "10010101100110",
                      23 when "10010101100111",
                      23 when "10010101101000",
                      23 when "10010101101001",
                      23 when "10010101101010",
                      23 when "10010101101011",
                      23 when "10010101101100",
                      23 when "10010101101101",
                      23 when "10010101101110",
                      23 when "10010101101111",
                      23 when "10010101110000",
                      23 when "10010101110001",
                      23 when "10010101110010",
                      23 when "10010101110011",
                      23 when "10010101110100",
                      23 when "10010101110101",
                      23 when "10010101110110",
                      23 when "10010101110111",
                      23 when "10010101111000",
                      23 when "10010101111001",
                      23 when "10010101111010",
                      23 when "10010101111011",
                      23 when "10010101111100",
                      23 when "10010101111101",
                      23 when "10010101111110",
                      23 when "10010101111111",
                      23 when "10010110000000",
                      23 when "10010110000001",
                      23 when "10010110000010",
                      23 when "10010110000011",
                      23 when "10010110000100",
                      23 when "10010110000101",
                      23 when "10010110000110",
                      23 when "10010110000111",
                      23 when "10010110001000",
                      23 when "10010110001001",
                      23 when "10010110001010",
                      23 when "10010110001011",
                      23 when "10010110001100",
                      23 when "10010110001101",
                      23 when "10010110001110",
                      23 when "10010110001111",
                      23 when "10010110010000",
                      23 when "10010110010001",
                      23 when "10010110010010",
                      23 when "10010110010011",
                      23 when "10010110010100",
                      23 when "10010110010101",
                      23 when "10010110010110",
                      23 when "10010110010111",
                      23 when "10010110011000",
                      23 when "10010110011001",
                      23 when "10010110011010",
                      23 when "10010110011011",
                      23 when "10010110011100",
                      23 when "10010110011101",
                      23 when "10010110011110",
                      23 when "10010110011111",
                      23 when "10010110100000",
                      23 when "10010110100001",
                      23 when "10010110100010",
                      23 when "10010110100011",
                      23 when "10010110100100",
                      23 when "10010110100101",
                      23 when "10010110100110",
                      23 when "10010110100111",
                      23 when "10010110101000",
                      23 when "10010110101001",
                      23 when "10010110101010",
                      23 when "10010110101011",
                      23 when "10010110101100",
                      23 when "10010110101101",
                      23 when "10010110101110",
                      23 when "10010110101111",
                      23 when "10010110110000",
                      23 when "10010110110001",
                      23 when "10010110110010",
                      23 when "10010110110011",
                      23 when "10010110110100",
                      23 when "10010110110101",
                      23 when "10010110110110",
                      23 when "10010110110111",
                      23 when "10010110111000",
                      23 when "10010110111001",
                      23 when "10010110111010",
                      23 when "10010110111011",
                      23 when "10010110111100",
                      23 when "10010110111101",
                      23 when "10010110111110",
                      23 when "10010110111111",
                      23 when "10010111000000",
                      23 when "10010111000001",
                      23 when "10010111000010",
                      23 when "10010111000011",
                      23 when "10010111000100",
                      23 when "10010111000101",
                      23 when "10010111000110",
                      23 when "10010111000111",
                      23 when "10010111001000",
                      23 when "10010111001001",
                      23 when "10010111001010",
                      23 when "10010111001011",
                      23 when "10010111001100",
                      23 when "10010111001101",
                      23 when "10010111001110",
                      23 when "10010111001111",
                      23 when "10010111010000",
                      23 when "10010111010001",
                      23 when "10010111010010",
                      23 when "10010111010011",
                      23 when "10010111010100",
                      23 when "10010111010101",
                      23 when "10010111010110",
                      23 when "10010111010111",
                      23 when "10010111011000",
                      23 when "10010111011001",
                      23 when "10010111011010",
                      23 when "10010111011011",
                      23 when "10010111011100",
                      23 when "10010111011101",
                      23 when "10010111011110",
                      23 when "10010111011111",
                      23 when "10010111100000",
                      23 when "10010111100001",
                      23 when "10010111100010",
                      23 when "10010111100011",
                      23 when "10010111100100",
                      23 when "10010111100101",
                      23 when "10010111100110",
                      23 when "10010111100111",
                      23 when "10010111101000",
                      23 when "10010111101001",
                      23 when "10010111101010",
                      23 when "10010111101011",
                      23 when "10010111101100",
                      23 when "10010111101101",
                      23 when "10010111101110",
                      23 when "10010111101111",
                      23 when "10010111110000",
                      23 when "10010111110001",
                      23 when "10010111110010",
                      23 when "10010111110011",
                      23 when "10010111110100",
                      23 when "10010111110101",
                      23 when "10010111110110",
                      23 when "10010111110111",
                      23 when "10010111111000",
                      23 when "10010111111001",
                      23 when "10010111111010",
                      23 when "10010111111011",
                      23 when "10010111111100",
                      23 when "10010111111101",
                      23 when "10010111111110",
                      23 when "10010111111111",
                      23 when "10011000000000",
                      23 when "10011000000001",
                      23 when "10011000000010",
                      23 when "10011000000011",
                      23 when "10011000000100",
                      23 when "10011000000101",
                      23 when "10011000000110",
                      23 when "10011000000111",
                      23 when "10011000001000",
                      23 when "10011000001001",
                      23 when "10011000001010",
                      23 when "10011000001011",
                      23 when "10011000001100",
                      23 when "10011000001101",
                      23 when "10011000001110",
                      23 when "10011000001111",
                      23 when "10011000010000",
                      23 when "10011000010001",
                      23 when "10011000010010",
                      23 when "10011000010011",
                      23 when "10011000010100",
                      23 when "10011000010101",
                      23 when "10011000010110",
                      23 when "10011000010111",
                      23 when "10011000011000",
                      23 when "10011000011001",
                      23 when "10011000011010",
                      23 when "10011000011011",
                      23 when "10011000011100",
                      23 when "10011000011101",
                      23 when "10011000011110",
                      23 when "10011000011111",
                      23 when "10011000100000",
                      23 when "10011000100001",
                      23 when "10011000100010",
                      23 when "10011000100011",
                      23 when "10011000100100",
                      23 when "10011000100101",
                      22 when "10011000100110",
                      22 when "10011000100111",
                      22 when "10011000101000",
                      22 when "10011000101001",
                      22 when "10011000101010",
                      22 when "10011000101011",
                      22 when "10011000101100",
                      22 when "10011000101101",
                      22 when "10011000101110",
                      22 when "10011000101111",
                      22 when "10011000110000",
                      22 when "10011000110001",
                      22 when "10011000110010",
                      22 when "10011000110011",
                      22 when "10011000110100",
                      22 when "10011000110101",
                      22 when "10011000110110",
                      22 when "10011000110111",
                      22 when "10011000111000",
                      22 when "10011000111001",
                      22 when "10011000111010",
                      22 when "10011000111011",
                      22 when "10011000111100",
                      22 when "10011000111101",
                      22 when "10011000111110",
                      22 when "10011000111111",
                      22 when "10011001000000",
                      22 when "10011001000001",
                      22 when "10011001000010",
                      22 when "10011001000011",
                      22 when "10011001000100",
                      22 when "10011001000101",
                      22 when "10011001000110",
                      22 when "10011001000111",
                      22 when "10011001001000",
                      22 when "10011001001001",
                      22 when "10011001001010",
                      22 when "10011001001011",
                      22 when "10011001001100",
                      22 when "10011001001101",
                      22 when "10011001001110",
                      22 when "10011001001111",
                      22 when "10011001010000",
                      22 when "10011001010001",
                      22 when "10011001010010",
                      22 when "10011001010011",
                      22 when "10011001010100",
                      22 when "10011001010101",
                      22 when "10011001010110",
                      22 when "10011001010111",
                      22 when "10011001011000",
                      22 when "10011001011001",
                      22 when "10011001011010",
                      22 when "10011001011011",
                      22 when "10011001011100",
                      22 when "10011001011101",
                      22 when "10011001011110",
                      22 when "10011001011111",
                      22 when "10011001100000",
                      22 when "10011001100001",
                      22 when "10011001100010",
                      22 when "10011001100011",
                      22 when "10011001100100",
                      22 when "10011001100101",
                      22 when "10011001100110",
                      22 when "10011001100111",
                      22 when "10011001101000",
                      22 when "10011001101001",
                      22 when "10011001101010",
                      22 when "10011001101011",
                      22 when "10011001101100",
                      22 when "10011001101101",
                      22 when "10011001101110",
                      22 when "10011001101111",
                      22 when "10011001110000",
                      22 when "10011001110001",
                      22 when "10011001110010",
                      22 when "10011001110011",
                      22 when "10011001110100",
                      22 when "10011001110101",
                      22 when "10011001110110",
                      22 when "10011001110111",
                      22 when "10011001111000",
                      22 when "10011001111001",
                      22 when "10011001111010",
                      22 when "10011001111011",
                      22 when "10011001111100",
                      22 when "10011001111101",
                      22 when "10011001111110",
                      22 when "10011001111111",
                      22 when "10011010000000",
                      22 when "10011010000001",
                      22 when "10011010000010",
                      22 when "10011010000011",
                      22 when "10011010000100",
                      22 when "10011010000101",
                      22 when "10011010000110",
                      22 when "10011010000111",
                      22 when "10011010001000",
                      22 when "10011010001001",
                      22 when "10011010001010",
                      22 when "10011010001011",
                      22 when "10011010001100",
                      22 when "10011010001101",
                      22 when "10011010001110",
                      22 when "10011010001111",
                      22 when "10011010010000",
                      22 when "10011010010001",
                      22 when "10011010010010",
                      22 when "10011010010011",
                      22 when "10011010010100",
                      22 when "10011010010101",
                      22 when "10011010010110",
                      22 when "10011010010111",
                      22 when "10011010011000",
                      22 when "10011010011001",
                      22 when "10011010011010",
                      22 when "10011010011011",
                      22 when "10011010011100",
                      22 when "10011010011101",
                      22 when "10011010011110",
                      22 when "10011010011111",
                      22 when "10011010100000",
                      22 when "10011010100001",
                      22 when "10011010100010",
                      22 when "10011010100011",
                      22 when "10011010100100",
                      22 when "10011010100101",
                      22 when "10011010100110",
                      22 when "10011010100111",
                      22 when "10011010101000",
                      22 when "10011010101001",
                      22 when "10011010101010",
                      22 when "10011010101011",
                      22 when "10011010101100",
                      22 when "10011010101101",
                      22 when "10011010101110",
                      22 when "10011010101111",
                      22 when "10011010110000",
                      22 when "10011010110001",
                      22 when "10011010110010",
                      22 when "10011010110011",
                      22 when "10011010110100",
                      22 when "10011010110101",
                      22 when "10011010110110",
                      22 when "10011010110111",
                      22 when "10011010111000",
                      22 when "10011010111001",
                      22 when "10011010111010",
                      22 when "10011010111011",
                      22 when "10011010111100",
                      22 when "10011010111101",
                      22 when "10011010111110",
                      22 when "10011010111111",
                      22 when "10011011000000",
                      22 when "10011011000001",
                      22 when "10011011000010",
                      22 when "10011011000011",
                      22 when "10011011000100",
                      22 when "10011011000101",
                      22 when "10011011000110",
                      22 when "10011011000111",
                      22 when "10011011001000",
                      22 when "10011011001001",
                      22 when "10011011001010",
                      22 when "10011011001011",
                      22 when "10011011001100",
                      22 when "10011011001101",
                      22 when "10011011001110",
                      22 when "10011011001111",
                      22 when "10011011010000",
                      22 when "10011011010001",
                      22 when "10011011010010",
                      22 when "10011011010011",
                      22 when "10011011010100",
                      22 when "10011011010101",
                      22 when "10011011010110",
                      22 when "10011011010111",
                      22 when "10011011011000",
                      22 when "10011011011001",
                      22 when "10011011011010",
                      22 when "10011011011011",
                      22 when "10011011011100",
                      22 when "10011011011101",
                      22 when "10011011011110",
                      22 when "10011011011111",
                      22 when "10011011100000",
                      22 when "10011011100001",
                      22 when "10011011100010",
                      22 when "10011011100011",
                      22 when "10011011100100",
                      22 when "10011011100101",
                      22 when "10011011100110",
                      22 when "10011011100111",
                      22 when "10011011101000",
                      22 when "10011011101001",
                      22 when "10011011101010",
                      22 when "10011011101011",
                      22 when "10011011101100",
                      22 when "10011011101101",
                      22 when "10011011101110",
                      22 when "10011011101111",
                      22 when "10011011110000",
                      22 when "10011011110001",
                      22 when "10011011110010",
                      22 when "10011011110011",
                      22 when "10011011110100",
                      22 when "10011011110101",
                      22 when "10011011110110",
                      22 when "10011011110111",
                      22 when "10011011111000",
                      22 when "10011011111001",
                      22 when "10011011111010",
                      22 when "10011011111011",
                      22 when "10011011111100",
                      22 when "10011011111101",
                      22 when "10011011111110",
                      22 when "10011011111111",
                      22 when "10011100000000",
                      22 when "10011100000001",
                      22 when "10011100000010",
                      22 when "10011100000011",
                      22 when "10011100000100",
                      22 when "10011100000101",
                      22 when "10011100000110",
                      22 when "10011100000111",
                      22 when "10011100001000",
                      22 when "10011100001001",
                      22 when "10011100001010",
                      22 when "10011100001011",
                      22 when "10011100001100",
                      22 when "10011100001101",
                      22 when "10011100001110",
                      22 when "10011100001111",
                      22 when "10011100010000",
                      22 when "10011100010001",
                      22 when "10011100010010",
                      22 when "10011100010011",
                      22 when "10011100010100",
                      22 when "10011100010101",
                      22 when "10011100010110",
                      22 when "10011100010111",
                      22 when "10011100011000",
                      22 when "10011100011001",
                      22 when "10011100011010",
                      22 when "10011100011011",
                      22 when "10011100011100",
                      22 when "10011100011101",
                      22 when "10011100011110",
                      22 when "10011100011111",
                      22 when "10011100100000",
                      22 when "10011100100001",
                      22 when "10011100100010",
                      22 when "10011100100011",
                      22 when "10011100100100",
                      22 when "10011100100101",
                      22 when "10011100100110",
                      22 when "10011100100111",
                      22 when "10011100101000",
                      22 when "10011100101001",
                      22 when "10011100101010",
                      22 when "10011100101011",
                      22 when "10011100101100",
                      22 when "10011100101101",
                      22 when "10011100101110",
                      22 when "10011100101111",
                      22 when "10011100110000",
                      22 when "10011100110001",
                      22 when "10011100110010",
                      22 when "10011100110011",
                      22 when "10011100110100",
                      22 when "10011100110101",
                      22 when "10011100110110",
                      22 when "10011100110111",
                      22 when "10011100111000",
                      22 when "10011100111001",
                      22 when "10011100111010",
                      22 when "10011100111011",
                      22 when "10011100111100",
                      22 when "10011100111101",
                      22 when "10011100111110",
                      22 when "10011100111111",
                      22 when "10011101000000",
                      22 when "10011101000001",
                      22 when "10011101000010",
                      22 when "10011101000011",
                      22 when "10011101000100",
                      22 when "10011101000101",
                      22 when "10011101000110",
                      22 when "10011101000111",
                      22 when "10011101001000",
                      22 when "10011101001001",
                      22 when "10011101001010",
                      22 when "10011101001011",
                      22 when "10011101001100",
                      22 when "10011101001101",
                      22 when "10011101001110",
                      22 when "10011101001111",
                      22 when "10011101010000",
                      22 when "10011101010001",
                      22 when "10011101010010",
                      22 when "10011101010011",
                      22 when "10011101010100",
                      22 when "10011101010101",
                      22 when "10011101010110",
                      22 when "10011101010111",
                      22 when "10011101011000",
                      22 when "10011101011001",
                      22 when "10011101011010",
                      22 when "10011101011011",
                      22 when "10011101011100",
                      22 when "10011101011101",
                      22 when "10011101011110",
                      22 when "10011101011111",
                      22 when "10011101100000",
                      22 when "10011101100001",
                      22 when "10011101100010",
                      22 when "10011101100011",
                      22 when "10011101100100",
                      22 when "10011101100101",
                      22 when "10011101100110",
                      22 when "10011101100111",
                      22 when "10011101101000",
                      22 when "10011101101001",
                      22 when "10011101101010",
                      22 when "10011101101011",
                      22 when "10011101101100",
                      22 when "10011101101101",
                      22 when "10011101101110",
                      22 when "10011101101111",
                      22 when "10011101110000",
                      22 when "10011101110001",
                      22 when "10011101110010",
                      22 when "10011101110011",
                      22 when "10011101110100",
                      22 when "10011101110101",
                      22 when "10011101110110",
                      22 when "10011101110111",
                      22 when "10011101111000",
                      22 when "10011101111001",
                      22 when "10011101111010",
                      22 when "10011101111011",
                      22 when "10011101111100",
                      22 when "10011101111101",
                      22 when "10011101111110",
                      22 when "10011101111111",
                      22 when "10011110000000",
                      22 when "10011110000001",
                      22 when "10011110000010",
                      22 when "10011110000011",
                      22 when "10011110000100",
                      22 when "10011110000101",
                      22 when "10011110000110",
                      22 when "10011110000111",
                      22 when "10011110001000",
                      22 when "10011110001001",
                      22 when "10011110001010",
                      22 when "10011110001011",
                      22 when "10011110001100",
                      22 when "10011110001101",
                      22 when "10011110001110",
                      22 when "10011110001111",
                      22 when "10011110010000",
                      22 when "10011110010001",
                      22 when "10011110010010",
                      22 when "10011110010011",
                      22 when "10011110010100",
                      22 when "10011110010101",
                      22 when "10011110010110",
                      22 when "10011110010111",
                      22 when "10011110011000",
                      22 when "10011110011001",
                      22 when "10011110011010",
                      22 when "10011110011011",
                      22 when "10011110011100",
                      22 when "10011110011101",
                      22 when "10011110011110",
                      22 when "10011110011111",
                      22 when "10011110100000",
                      22 when "10011110100001",
                      22 when "10011110100010",
                      22 when "10011110100011",
                      22 when "10011110100100",
                      22 when "10011110100101",
                      22 when "10011110100110",
                      22 when "10011110100111",
                      22 when "10011110101000",
                      22 when "10011110101001",
                      22 when "10011110101010",
                      22 when "10011110101011",
                      22 when "10011110101100",
                      22 when "10011110101101",
                      22 when "10011110101110",
                      22 when "10011110101111",
                      22 when "10011110110000",
                      22 when "10011110110001",
                      22 when "10011110110010",
                      22 when "10011110110011",
                      22 when "10011110110100",
                      22 when "10011110110101",
                      22 when "10011110110110",
                      22 when "10011110110111",
                      22 when "10011110111000",
                      22 when "10011110111001",
                      22 when "10011110111010",
                      22 when "10011110111011",
                      22 when "10011110111100",
                      22 when "10011110111101",
                      22 when "10011110111110",
                      22 when "10011110111111",
                      22 when "10011111000000",
                      22 when "10011111000001",
                      22 when "10011111000010",
                      22 when "10011111000011",
                      22 when "10011111000100",
                      22 when "10011111000101",
                      22 when "10011111000110",
                      22 when "10011111000111",
                      22 when "10011111001000",
                      22 when "10011111001001",
                      22 when "10011111001010",
                      22 when "10011111001011",
                      22 when "10011111001100",
                      22 when "10011111001101",
                      22 when "10011111001110",
                      22 when "10011111001111",
                      22 when "10011111010000",
                      22 when "10011111010001",
                      22 when "10011111010010",
                      22 when "10011111010011",
                      22 when "10011111010100",
                      22 when "10011111010101",
                      22 when "10011111010110",
                      22 when "10011111010111",
                      22 when "10011111011000",
                      22 when "10011111011001",
                      22 when "10011111011010",
                      22 when "10011111011011",
                      22 when "10011111011100",
                      22 when "10011111011101",
                      22 when "10011111011110",
                      22 when "10011111011111",
                      22 when "10011111100000",
                      22 when "10011111100001",
                      22 when "10011111100010",
                      22 when "10011111100011",
                      22 when "10011111100100",
                      22 when "10011111100101",
                      22 when "10011111100110",
                      22 when "10011111100111",
                      22 when "10011111101000",
                      22 when "10011111101001",
                      22 when "10011111101010",
                      22 when "10011111101011",
                      21 when "10011111101100",
                      21 when "10011111101101",
                      21 when "10011111101110",
                      21 when "10011111101111",
                      21 when "10011111110000",
                      21 when "10011111110001",
                      21 when "10011111110010",
                      21 when "10011111110011",
                      21 when "10011111110100",
                      21 when "10011111110101",
                      21 when "10011111110110",
                      21 when "10011111110111",
                      21 when "10011111111000",
                      21 when "10011111111001",
                      21 when "10011111111010",
                      21 when "10011111111011",
                      21 when "10011111111100",
                      21 when "10011111111101",
                      21 when "10011111111110",
                      21 when "10011111111111",
                      21 when "10100000000000",
                      21 when "10100000000001",
                      21 when "10100000000010",
                      21 when "10100000000011",
                      21 when "10100000000100",
                      21 when "10100000000101",
                      21 when "10100000000110",
                      21 when "10100000000111",
                      21 when "10100000001000",
                      21 when "10100000001001",
                      21 when "10100000001010",
                      21 when "10100000001011",
                      21 when "10100000001100",
                      21 when "10100000001101",
                      21 when "10100000001110",
                      21 when "10100000001111",
                      21 when "10100000010000",
                      21 when "10100000010001",
                      21 when "10100000010010",
                      21 when "10100000010011",
                      21 when "10100000010100",
                      21 when "10100000010101",
                      21 when "10100000010110",
                      21 when "10100000010111",
                      21 when "10100000011000",
                      21 when "10100000011001",
                      21 when "10100000011010",
                      21 when "10100000011011",
                      21 when "10100000011100",
                      21 when "10100000011101",
                      21 when "10100000011110",
                      21 when "10100000011111",
                      21 when "10100000100000",
                      21 when "10100000100001",
                      21 when "10100000100010",
                      21 when "10100000100011",
                      21 when "10100000100100",
                      21 when "10100000100101",
                      21 when "10100000100110",
                      21 when "10100000100111",
                      21 when "10100000101000",
                      21 when "10100000101001",
                      21 when "10100000101010",
                      21 when "10100000101011",
                      21 when "10100000101100",
                      21 when "10100000101101",
                      21 when "10100000101110",
                      21 when "10100000101111",
                      21 when "10100000110000",
                      21 when "10100000110001",
                      21 when "10100000110010",
                      21 when "10100000110011",
                      21 when "10100000110100",
                      21 when "10100000110101",
                      21 when "10100000110110",
                      21 when "10100000110111",
                      21 when "10100000111000",
                      21 when "10100000111001",
                      21 when "10100000111010",
                      21 when "10100000111011",
                      21 when "10100000111100",
                      21 when "10100000111101",
                      21 when "10100000111110",
                      21 when "10100000111111",
                      21 when "10100001000000",
                      21 when "10100001000001",
                      21 when "10100001000010",
                      21 when "10100001000011",
                      21 when "10100001000100",
                      21 when "10100001000101",
                      21 when "10100001000110",
                      21 when "10100001000111",
                      21 when "10100001001000",
                      21 when "10100001001001",
                      21 when "10100001001010",
                      21 when "10100001001011",
                      21 when "10100001001100",
                      21 when "10100001001101",
                      21 when "10100001001110",
                      21 when "10100001001111",
                      21 when "10100001010000",
                      21 when "10100001010001",
                      21 when "10100001010010",
                      21 when "10100001010011",
                      21 when "10100001010100",
                      21 when "10100001010101",
                      21 when "10100001010110",
                      21 when "10100001010111",
                      21 when "10100001011000",
                      21 when "10100001011001",
                      21 when "10100001011010",
                      21 when "10100001011011",
                      21 when "10100001011100",
                      21 when "10100001011101",
                      21 when "10100001011110",
                      21 when "10100001011111",
                      21 when "10100001100000",
                      21 when "10100001100001",
                      21 when "10100001100010",
                      21 when "10100001100011",
                      21 when "10100001100100",
                      21 when "10100001100101",
                      21 when "10100001100110",
                      21 when "10100001100111",
                      21 when "10100001101000",
                      21 when "10100001101001",
                      21 when "10100001101010",
                      21 when "10100001101011",
                      21 when "10100001101100",
                      21 when "10100001101101",
                      21 when "10100001101110",
                      21 when "10100001101111",
                      21 when "10100001110000",
                      21 when "10100001110001",
                      21 when "10100001110010",
                      21 when "10100001110011",
                      21 when "10100001110100",
                      21 when "10100001110101",
                      21 when "10100001110110",
                      21 when "10100001110111",
                      21 when "10100001111000",
                      21 when "10100001111001",
                      21 when "10100001111010",
                      21 when "10100001111011",
                      21 when "10100001111100",
                      21 when "10100001111101",
                      21 when "10100001111110",
                      21 when "10100001111111",
                      21 when "10100010000000",
                      21 when "10100010000001",
                      21 when "10100010000010",
                      21 when "10100010000011",
                      21 when "10100010000100",
                      21 when "10100010000101",
                      21 when "10100010000110",
                      21 when "10100010000111",
                      21 when "10100010001000",
                      21 when "10100010001001",
                      21 when "10100010001010",
                      21 when "10100010001011",
                      21 when "10100010001100",
                      21 when "10100010001101",
                      21 when "10100010001110",
                      21 when "10100010001111",
                      21 when "10100010010000",
                      21 when "10100010010001",
                      21 when "10100010010010",
                      21 when "10100010010011",
                      21 when "10100010010100",
                      21 when "10100010010101",
                      21 when "10100010010110",
                      21 when "10100010010111",
                      21 when "10100010011000",
                      21 when "10100010011001",
                      21 when "10100010011010",
                      21 when "10100010011011",
                      21 when "10100010011100",
                      21 when "10100010011101",
                      21 when "10100010011110",
                      21 when "10100010011111",
                      21 when "10100010100000",
                      21 when "10100010100001",
                      21 when "10100010100010",
                      21 when "10100010100011",
                      21 when "10100010100100",
                      21 when "10100010100101",
                      21 when "10100010100110",
                      21 when "10100010100111",
                      21 when "10100010101000",
                      21 when "10100010101001",
                      21 when "10100010101010",
                      21 when "10100010101011",
                      21 when "10100010101100",
                      21 when "10100010101101",
                      21 when "10100010101110",
                      21 when "10100010101111",
                      21 when "10100010110000",
                      21 when "10100010110001",
                      21 when "10100010110010",
                      21 when "10100010110011",
                      21 when "10100010110100",
                      21 when "10100010110101",
                      21 when "10100010110110",
                      21 when "10100010110111",
                      21 when "10100010111000",
                      21 when "10100010111001",
                      21 when "10100010111010",
                      21 when "10100010111011",
                      21 when "10100010111100",
                      21 when "10100010111101",
                      21 when "10100010111110",
                      21 when "10100010111111",
                      21 when "10100011000000",
                      21 when "10100011000001",
                      21 when "10100011000010",
                      21 when "10100011000011",
                      21 when "10100011000100",
                      21 when "10100011000101",
                      21 when "10100011000110",
                      21 when "10100011000111",
                      21 when "10100011001000",
                      21 when "10100011001001",
                      21 when "10100011001010",
                      21 when "10100011001011",
                      21 when "10100011001100",
                      21 when "10100011001101",
                      21 when "10100011001110",
                      21 when "10100011001111",
                      21 when "10100011010000",
                      21 when "10100011010001",
                      21 when "10100011010010",
                      21 when "10100011010011",
                      21 when "10100011010100",
                      21 when "10100011010101",
                      21 when "10100011010110",
                      21 when "10100011010111",
                      21 when "10100011011000",
                      21 when "10100011011001",
                      21 when "10100011011010",
                      21 when "10100011011011",
                      21 when "10100011011100",
                      21 when "10100011011101",
                      21 when "10100011011110",
                      21 when "10100011011111",
                      21 when "10100011100000",
                      21 when "10100011100001",
                      21 when "10100011100010",
                      21 when "10100011100011",
                      21 when "10100011100100",
                      21 when "10100011100101",
                      21 when "10100011100110",
                      21 when "10100011100111",
                      21 when "10100011101000",
                      21 when "10100011101001",
                      21 when "10100011101010",
                      21 when "10100011101011",
                      21 when "10100011101100",
                      21 when "10100011101101",
                      21 when "10100011101110",
                      21 when "10100011101111",
                      21 when "10100011110000",
                      21 when "10100011110001",
                      21 when "10100011110010",
                      21 when "10100011110011",
                      21 when "10100011110100",
                      21 when "10100011110101",
                      21 when "10100011110110",
                      21 when "10100011110111",
                      21 when "10100011111000",
                      21 when "10100011111001",
                      21 when "10100011111010",
                      21 when "10100011111011",
                      21 when "10100011111100",
                      21 when "10100011111101",
                      21 when "10100011111110",
                      21 when "10100011111111",
                      21 when "10100100000000",
                      21 when "10100100000001",
                      21 when "10100100000010",
                      21 when "10100100000011",
                      21 when "10100100000100",
                      21 when "10100100000101",
                      21 when "10100100000110",
                      21 when "10100100000111",
                      21 when "10100100001000",
                      21 when "10100100001001",
                      21 when "10100100001010",
                      21 when "10100100001011",
                      21 when "10100100001100",
                      21 when "10100100001101",
                      21 when "10100100001110",
                      21 when "10100100001111",
                      21 when "10100100010000",
                      21 when "10100100010001",
                      21 when "10100100010010",
                      21 when "10100100010011",
                      21 when "10100100010100",
                      21 when "10100100010101",
                      21 when "10100100010110",
                      21 when "10100100010111",
                      21 when "10100100011000",
                      21 when "10100100011001",
                      21 when "10100100011010",
                      21 when "10100100011011",
                      21 when "10100100011100",
                      21 when "10100100011101",
                      21 when "10100100011110",
                      21 when "10100100011111",
                      21 when "10100100100000",
                      21 when "10100100100001",
                      21 when "10100100100010",
                      21 when "10100100100011",
                      21 when "10100100100100",
                      21 when "10100100100101",
                      21 when "10100100100110",
                      21 when "10100100100111",
                      21 when "10100100101000",
                      21 when "10100100101001",
                      21 when "10100100101010",
                      21 when "10100100101011",
                      21 when "10100100101100",
                      21 when "10100100101101",
                      21 when "10100100101110",
                      21 when "10100100101111",
                      21 when "10100100110000",
                      21 when "10100100110001",
                      21 when "10100100110010",
                      21 when "10100100110011",
                      21 when "10100100110100",
                      21 when "10100100110101",
                      21 when "10100100110110",
                      21 when "10100100110111",
                      21 when "10100100111000",
                      21 when "10100100111001",
                      21 when "10100100111010",
                      21 when "10100100111011",
                      21 when "10100100111100",
                      21 when "10100100111101",
                      21 when "10100100111110",
                      21 when "10100100111111",
                      21 when "10100101000000",
                      21 when "10100101000001",
                      21 when "10100101000010",
                      21 when "10100101000011",
                      21 when "10100101000100",
                      21 when "10100101000101",
                      21 when "10100101000110",
                      21 when "10100101000111",
                      21 when "10100101001000",
                      21 when "10100101001001",
                      21 when "10100101001010",
                      21 when "10100101001011",
                      21 when "10100101001100",
                      21 when "10100101001101",
                      21 when "10100101001110",
                      21 when "10100101001111",
                      21 when "10100101010000",
                      21 when "10100101010001",
                      21 when "10100101010010",
                      21 when "10100101010011",
                      21 when "10100101010100",
                      21 when "10100101010101",
                      21 when "10100101010110",
                      21 when "10100101010111",
                      21 when "10100101011000",
                      21 when "10100101011001",
                      21 when "10100101011010",
                      21 when "10100101011011",
                      21 when "10100101011100",
                      21 when "10100101011101",
                      21 when "10100101011110",
                      21 when "10100101011111",
                      21 when "10100101100000",
                      21 when "10100101100001",
                      21 when "10100101100010",
                      21 when "10100101100011",
                      21 when "10100101100100",
                      21 when "10100101100101",
                      21 when "10100101100110",
                      21 when "10100101100111",
                      21 when "10100101101000",
                      21 when "10100101101001",
                      21 when "10100101101010",
                      21 when "10100101101011",
                      21 when "10100101101100",
                      21 when "10100101101101",
                      21 when "10100101101110",
                      21 when "10100101101111",
                      21 when "10100101110000",
                      21 when "10100101110001",
                      21 when "10100101110010",
                      21 when "10100101110011",
                      21 when "10100101110100",
                      21 when "10100101110101",
                      21 when "10100101110110",
                      21 when "10100101110111",
                      21 when "10100101111000",
                      21 when "10100101111001",
                      21 when "10100101111010",
                      21 when "10100101111011",
                      21 when "10100101111100",
                      21 when "10100101111101",
                      21 when "10100101111110",
                      21 when "10100101111111",
                      21 when "10100110000000",
                      21 when "10100110000001",
                      21 when "10100110000010",
                      21 when "10100110000011",
                      21 when "10100110000100",
                      21 when "10100110000101",
                      21 when "10100110000110",
                      21 when "10100110000111",
                      21 when "10100110001000",
                      21 when "10100110001001",
                      21 when "10100110001010",
                      21 when "10100110001011",
                      21 when "10100110001100",
                      21 when "10100110001101",
                      21 when "10100110001110",
                      21 when "10100110001111",
                      21 when "10100110010000",
                      21 when "10100110010001",
                      21 when "10100110010010",
                      21 when "10100110010011",
                      21 when "10100110010100",
                      21 when "10100110010101",
                      21 when "10100110010110",
                      21 when "10100110010111",
                      21 when "10100110011000",
                      21 when "10100110011001",
                      21 when "10100110011010",
                      21 when "10100110011011",
                      21 when "10100110011100",
                      21 when "10100110011101",
                      21 when "10100110011110",
                      21 when "10100110011111",
                      21 when "10100110100000",
                      21 when "10100110100001",
                      21 when "10100110100010",
                      21 when "10100110100011",
                      21 when "10100110100100",
                      21 when "10100110100101",
                      21 when "10100110100110",
                      21 when "10100110100111",
                      21 when "10100110101000",
                      21 when "10100110101001",
                      21 when "10100110101010",
                      21 when "10100110101011",
                      21 when "10100110101100",
                      21 when "10100110101101",
                      21 when "10100110101110",
                      21 when "10100110101111",
                      21 when "10100110110000",
                      21 when "10100110110001",
                      21 when "10100110110010",
                      21 when "10100110110011",
                      21 when "10100110110100",
                      21 when "10100110110101",
                      21 when "10100110110110",
                      21 when "10100110110111",
                      21 when "10100110111000",
                      21 when "10100110111001",
                      21 when "10100110111010",
                      21 when "10100110111011",
                      21 when "10100110111100",
                      21 when "10100110111101",
                      21 when "10100110111110",
                      21 when "10100110111111",
                      21 when "10100111000000",
                      21 when "10100111000001",
                      21 when "10100111000010",
                      21 when "10100111000011",
                      21 when "10100111000100",
                      21 when "10100111000101",
                      21 when "10100111000110",
                      21 when "10100111000111",
                      21 when "10100111001000",
                      21 when "10100111001001",
                      21 when "10100111001010",
                      21 when "10100111001011",
                      21 when "10100111001100",
                      21 when "10100111001101",
                      21 when "10100111001110",
                      21 when "10100111001111",
                      21 when "10100111010000",
                      21 when "10100111010001",
                      21 when "10100111010010",
                      21 when "10100111010011",
                      21 when "10100111010100",
                      21 when "10100111010101",
                      21 when "10100111010110",
                      21 when "10100111010111",
                      21 when "10100111011000",
                      21 when "10100111011001",
                      21 when "10100111011010",
                      21 when "10100111011011",
                      21 when "10100111011100",
                      21 when "10100111011101",
                      21 when "10100111011110",
                      20 when "10100111011111",
                      20 when "10100111100000",
                      20 when "10100111100001",
                      20 when "10100111100010",
                      20 when "10100111100011",
                      20 when "10100111100100",
                      20 when "10100111100101",
                      20 when "10100111100110",
                      20 when "10100111100111",
                      20 when "10100111101000",
                      20 when "10100111101001",
                      20 when "10100111101010",
                      20 when "10100111101011",
                      20 when "10100111101100",
                      20 when "10100111101101",
                      20 when "10100111101110",
                      20 when "10100111101111",
                      20 when "10100111110000",
                      20 when "10100111110001",
                      20 when "10100111110010",
                      20 when "10100111110011",
                      20 when "10100111110100",
                      20 when "10100111110101",
                      20 when "10100111110110",
                      20 when "10100111110111",
                      20 when "10100111111000",
                      20 when "10100111111001",
                      20 when "10100111111010",
                      20 when "10100111111011",
                      20 when "10100111111100",
                      20 when "10100111111101",
                      20 when "10100111111110",
                      20 when "10100111111111",
                      20 when "10101000000000",
                      20 when "10101000000001",
                      20 when "10101000000010",
                      20 when "10101000000011",
                      20 when "10101000000100",
                      20 when "10101000000101",
                      20 when "10101000000110",
                      20 when "10101000000111",
                      20 when "10101000001000",
                      20 when "10101000001001",
                      20 when "10101000001010",
                      20 when "10101000001011",
                      20 when "10101000001100",
                      20 when "10101000001101",
                      20 when "10101000001110",
                      20 when "10101000001111",
                      20 when "10101000010000",
                      20 when "10101000010001",
                      20 when "10101000010010",
                      20 when "10101000010011",
                      20 when "10101000010100",
                      20 when "10101000010101",
                      20 when "10101000010110",
                      20 when "10101000010111",
                      20 when "10101000011000",
                      20 when "10101000011001",
                      20 when "10101000011010",
                      20 when "10101000011011",
                      20 when "10101000011100",
                      20 when "10101000011101",
                      20 when "10101000011110",
                      20 when "10101000011111",
                      20 when "10101000100000",
                      20 when "10101000100001",
                      20 when "10101000100010",
                      20 when "10101000100011",
                      20 when "10101000100100",
                      20 when "10101000100101",
                      20 when "10101000100110",
                      20 when "10101000100111",
                      20 when "10101000101000",
                      20 when "10101000101001",
                      20 when "10101000101010",
                      20 when "10101000101011",
                      20 when "10101000101100",
                      20 when "10101000101101",
                      20 when "10101000101110",
                      20 when "10101000101111",
                      20 when "10101000110000",
                      20 when "10101000110001",
                      20 when "10101000110010",
                      20 when "10101000110011",
                      20 when "10101000110100",
                      20 when "10101000110101",
                      20 when "10101000110110",
                      20 when "10101000110111",
                      20 when "10101000111000",
                      20 when "10101000111001",
                      20 when "10101000111010",
                      20 when "10101000111011",
                      20 when "10101000111100",
                      20 when "10101000111101",
                      20 when "10101000111110",
                      20 when "10101000111111",
                      20 when "10101001000000",
                      20 when "10101001000001",
                      20 when "10101001000010",
                      20 when "10101001000011",
                      20 when "10101001000100",
                      20 when "10101001000101",
                      20 when "10101001000110",
                      20 when "10101001000111",
                      20 when "10101001001000",
                      20 when "10101001001001",
                      20 when "10101001001010",
                      20 when "10101001001011",
                      20 when "10101001001100",
                      20 when "10101001001101",
                      20 when "10101001001110",
                      20 when "10101001001111",
                      20 when "10101001010000",
                      20 when "10101001010001",
                      20 when "10101001010010",
                      20 when "10101001010011",
                      20 when "10101001010100",
                      20 when "10101001010101",
                      20 when "10101001010110",
                      20 when "10101001010111",
                      20 when "10101001011000",
                      20 when "10101001011001",
                      20 when "10101001011010",
                      20 when "10101001011011",
                      20 when "10101001011100",
                      20 when "10101001011101",
                      20 when "10101001011110",
                      20 when "10101001011111",
                      20 when "10101001100000",
                      20 when "10101001100001",
                      20 when "10101001100010",
                      20 when "10101001100011",
                      20 when "10101001100100",
                      20 when "10101001100101",
                      20 when "10101001100110",
                      20 when "10101001100111",
                      20 when "10101001101000",
                      20 when "10101001101001",
                      20 when "10101001101010",
                      20 when "10101001101011",
                      20 when "10101001101100",
                      20 when "10101001101101",
                      20 when "10101001101110",
                      20 when "10101001101111",
                      20 when "10101001110000",
                      20 when "10101001110001",
                      20 when "10101001110010",
                      20 when "10101001110011",
                      20 when "10101001110100",
                      20 when "10101001110101",
                      20 when "10101001110110",
                      20 when "10101001110111",
                      20 when "10101001111000",
                      20 when "10101001111001",
                      20 when "10101001111010",
                      20 when "10101001111011",
                      20 when "10101001111100",
                      20 when "10101001111101",
                      20 when "10101001111110",
                      20 when "10101001111111",
                      20 when "10101010000000",
                      20 when "10101010000001",
                      20 when "10101010000010",
                      20 when "10101010000011",
                      20 when "10101010000100",
                      20 when "10101010000101",
                      20 when "10101010000110",
                      20 when "10101010000111",
                      20 when "10101010001000",
                      20 when "10101010001001",
                      20 when "10101010001010",
                      20 when "10101010001011",
                      20 when "10101010001100",
                      20 when "10101010001101",
                      20 when "10101010001110",
                      20 when "10101010001111",
                      20 when "10101010010000",
                      20 when "10101010010001",
                      20 when "10101010010010",
                      20 when "10101010010011",
                      20 when "10101010010100",
                      20 when "10101010010101",
                      20 when "10101010010110",
                      20 when "10101010010111",
                      20 when "10101010011000",
                      20 when "10101010011001",
                      20 when "10101010011010",
                      20 when "10101010011011",
                      20 when "10101010011100",
                      20 when "10101010011101",
                      20 when "10101010011110",
                      20 when "10101010011111",
                      20 when "10101010100000",
                      20 when "10101010100001",
                      20 when "10101010100010",
                      20 when "10101010100011",
                      20 when "10101010100100",
                      20 when "10101010100101",
                      20 when "10101010100110",
                      20 when "10101010100111",
                      20 when "10101010101000",
                      20 when "10101010101001",
                      20 when "10101010101010",
                      20 when "10101010101011",
                      20 when "10101010101100",
                      20 when "10101010101101",
                      20 when "10101010101110",
                      20 when "10101010101111",
                      20 when "10101010110000",
                      20 when "10101010110001",
                      20 when "10101010110010",
                      20 when "10101010110011",
                      20 when "10101010110100",
                      20 when "10101010110101",
                      20 when "10101010110110",
                      20 when "10101010110111",
                      20 when "10101010111000",
                      20 when "10101010111001",
                      20 when "10101010111010",
                      20 when "10101010111011",
                      20 when "10101010111100",
                      20 when "10101010111101",
                      20 when "10101010111110",
                      20 when "10101010111111",
                      20 when "10101011000000",
                      20 when "10101011000001",
                      20 when "10101011000010",
                      20 when "10101011000011",
                      20 when "10101011000100",
                      20 when "10101011000101",
                      20 when "10101011000110",
                      20 when "10101011000111",
                      20 when "10101011001000",
                      20 when "10101011001001",
                      20 when "10101011001010",
                      20 when "10101011001011",
                      20 when "10101011001100",
                      20 when "10101011001101",
                      20 when "10101011001110",
                      20 when "10101011001111",
                      20 when "10101011010000",
                      20 when "10101011010001",
                      20 when "10101011010010",
                      20 when "10101011010011",
                      20 when "10101011010100",
                      20 when "10101011010101",
                      20 when "10101011010110",
                      20 when "10101011010111",
                      20 when "10101011011000",
                      20 when "10101011011001",
                      20 when "10101011011010",
                      20 when "10101011011011",
                      20 when "10101011011100",
                      20 when "10101011011101",
                      20 when "10101011011110",
                      20 when "10101011011111",
                      20 when "10101011100000",
                      20 when "10101011100001",
                      20 when "10101011100010",
                      20 when "10101011100011",
                      20 when "10101011100100",
                      20 when "10101011100101",
                      20 when "10101011100110",
                      20 when "10101011100111",
                      20 when "10101011101000",
                      20 when "10101011101001",
                      20 when "10101011101010",
                      20 when "10101011101011",
                      20 when "10101011101100",
                      20 when "10101011101101",
                      20 when "10101011101110",
                      20 when "10101011101111",
                      20 when "10101011110000",
                      20 when "10101011110001",
                      20 when "10101011110010",
                      20 when "10101011110011",
                      20 when "10101011110100",
                      20 when "10101011110101",
                      20 when "10101011110110",
                      20 when "10101011110111",
                      20 when "10101011111000",
                      20 when "10101011111001",
                      20 when "10101011111010",
                      20 when "10101011111011",
                      20 when "10101011111100",
                      20 when "10101011111101",
                      20 when "10101011111110",
                      20 when "10101011111111",
                      20 when "10101100000000",
                      20 when "10101100000001",
                      20 when "10101100000010",
                      20 when "10101100000011",
                      20 when "10101100000100",
                      20 when "10101100000101",
                      20 when "10101100000110",
                      20 when "10101100000111",
                      20 when "10101100001000",
                      20 when "10101100001001",
                      20 when "10101100001010",
                      20 when "10101100001011",
                      20 when "10101100001100",
                      20 when "10101100001101",
                      20 when "10101100001110",
                      20 when "10101100001111",
                      20 when "10101100010000",
                      20 when "10101100010001",
                      20 when "10101100010010",
                      20 when "10101100010011",
                      20 when "10101100010100",
                      20 when "10101100010101",
                      20 when "10101100010110",
                      20 when "10101100010111",
                      20 when "10101100011000",
                      20 when "10101100011001",
                      20 when "10101100011010",
                      20 when "10101100011011",
                      20 when "10101100011100",
                      20 when "10101100011101",
                      20 when "10101100011110",
                      20 when "10101100011111",
                      20 when "10101100100000",
                      20 when "10101100100001",
                      20 when "10101100100010",
                      20 when "10101100100011",
                      20 when "10101100100100",
                      20 when "10101100100101",
                      20 when "10101100100110",
                      20 when "10101100100111",
                      20 when "10101100101000",
                      20 when "10101100101001",
                      20 when "10101100101010",
                      20 when "10101100101011",
                      20 when "10101100101100",
                      20 when "10101100101101",
                      20 when "10101100101110",
                      20 when "10101100101111",
                      20 when "10101100110000",
                      20 when "10101100110001",
                      20 when "10101100110010",
                      20 when "10101100110011",
                      20 when "10101100110100",
                      20 when "10101100110101",
                      20 when "10101100110110",
                      20 when "10101100110111",
                      20 when "10101100111000",
                      20 when "10101100111001",
                      20 when "10101100111010",
                      20 when "10101100111011",
                      20 when "10101100111100",
                      20 when "10101100111101",
                      20 when "10101100111110",
                      20 when "10101100111111",
                      20 when "10101101000000",
                      20 when "10101101000001",
                      20 when "10101101000010",
                      20 when "10101101000011",
                      20 when "10101101000100",
                      20 when "10101101000101",
                      20 when "10101101000110",
                      20 when "10101101000111",
                      20 when "10101101001000",
                      20 when "10101101001001",
                      20 when "10101101001010",
                      20 when "10101101001011",
                      20 when "10101101001100",
                      20 when "10101101001101",
                      20 when "10101101001110",
                      20 when "10101101001111",
                      20 when "10101101010000",
                      20 when "10101101010001",
                      20 when "10101101010010",
                      20 when "10101101010011",
                      20 when "10101101010100",
                      20 when "10101101010101",
                      20 when "10101101010110",
                      20 when "10101101010111",
                      20 when "10101101011000",
                      20 when "10101101011001",
                      20 when "10101101011010",
                      20 when "10101101011011",
                      20 when "10101101011100",
                      20 when "10101101011101",
                      20 when "10101101011110",
                      20 when "10101101011111",
                      20 when "10101101100000",
                      20 when "10101101100001",
                      20 when "10101101100010",
                      20 when "10101101100011",
                      20 when "10101101100100",
                      20 when "10101101100101",
                      20 when "10101101100110",
                      20 when "10101101100111",
                      20 when "10101101101000",
                      20 when "10101101101001",
                      20 when "10101101101010",
                      20 when "10101101101011",
                      20 when "10101101101100",
                      20 when "10101101101101",
                      20 when "10101101101110",
                      20 when "10101101101111",
                      20 when "10101101110000",
                      20 when "10101101110001",
                      20 when "10101101110010",
                      20 when "10101101110011",
                      20 when "10101101110100",
                      20 when "10101101110101",
                      20 when "10101101110110",
                      20 when "10101101110111",
                      20 when "10101101111000",
                      20 when "10101101111001",
                      20 when "10101101111010",
                      20 when "10101101111011",
                      20 when "10101101111100",
                      20 when "10101101111101",
                      20 when "10101101111110",
                      20 when "10101101111111",
                      20 when "10101110000000",
                      20 when "10101110000001",
                      20 when "10101110000010",
                      20 when "10101110000011",
                      20 when "10101110000100",
                      20 when "10101110000101",
                      20 when "10101110000110",
                      20 when "10101110000111",
                      20 when "10101110001000",
                      20 when "10101110001001",
                      20 when "10101110001010",
                      20 when "10101110001011",
                      20 when "10101110001100",
                      20 when "10101110001101",
                      20 when "10101110001110",
                      20 when "10101110001111",
                      20 when "10101110010000",
                      20 when "10101110010001",
                      20 when "10101110010010",
                      20 when "10101110010011",
                      20 when "10101110010100",
                      20 when "10101110010101",
                      20 when "10101110010110",
                      20 when "10101110010111",
                      20 when "10101110011000",
                      20 when "10101110011001",
                      20 when "10101110011010",
                      20 when "10101110011011",
                      20 when "10101110011100",
                      20 when "10101110011101",
                      20 when "10101110011110",
                      20 when "10101110011111",
                      20 when "10101110100000",
                      20 when "10101110100001",
                      20 when "10101110100010",
                      20 when "10101110100011",
                      20 when "10101110100100",
                      20 when "10101110100101",
                      20 when "10101110100110",
                      20 when "10101110100111",
                      20 when "10101110101000",
                      20 when "10101110101001",
                      20 when "10101110101010",
                      20 when "10101110101011",
                      20 when "10101110101100",
                      20 when "10101110101101",
                      20 when "10101110101110",
                      20 when "10101110101111",
                      20 when "10101110110000",
                      20 when "10101110110001",
                      20 when "10101110110010",
                      20 when "10101110110011",
                      20 when "10101110110100",
                      20 when "10101110110101",
                      20 when "10101110110110",
                      20 when "10101110110111",
                      20 when "10101110111000",
                      20 when "10101110111001",
                      20 when "10101110111010",
                      20 when "10101110111011",
                      20 when "10101110111100",
                      20 when "10101110111101",
                      20 when "10101110111110",
                      20 when "10101110111111",
                      20 when "10101111000000",
                      20 when "10101111000001",
                      20 when "10101111000010",
                      20 when "10101111000011",
                      20 when "10101111000100",
                      20 when "10101111000101",
                      20 when "10101111000110",
                      20 when "10101111000111",
                      20 when "10101111001000",
                      20 when "10101111001001",
                      20 when "10101111001010",
                      20 when "10101111001011",
                      20 when "10101111001100",
                      20 when "10101111001101",
                      20 when "10101111001110",
                      20 when "10101111001111",
                      20 when "10101111010000",
                      20 when "10101111010001",
                      20 when "10101111010010",
                      20 when "10101111010011",
                      20 when "10101111010100",
                      20 when "10101111010101",
                      20 when "10101111010110",
                      20 when "10101111010111",
                      20 when "10101111011000",
                      20 when "10101111011001",
                      20 when "10101111011010",
                      20 when "10101111011011",
                      20 when "10101111011100",
                      20 when "10101111011101",
                      20 when "10101111011110",
                      20 when "10101111011111",
                      20 when "10101111100000",
                      20 when "10101111100001",
                      20 when "10101111100010",
                      20 when "10101111100011",
                      20 when "10101111100100",
                      20 when "10101111100101",
                      20 when "10101111100110",
                      20 when "10101111100111",
                      20 when "10101111101000",
                      20 when "10101111101001",
                      20 when "10101111101010",
                      20 when "10101111101011",
                      20 when "10101111101100",
                      20 when "10101111101101",
                      20 when "10101111101110",
                      20 when "10101111101111",
                      20 when "10101111110000",
                      20 when "10101111110001",
                      20 when "10101111110010",
                      20 when "10101111110011",
                      20 when "10101111110100",
                      20 when "10101111110101",
                      20 when "10101111110110",
                      20 when "10101111110111",
                      20 when "10101111111000",
                      20 when "10101111111001",
                      20 when "10101111111010",
                      20 when "10101111111011",
                      20 when "10101111111100",
                      20 when "10101111111101",
                      20 when "10101111111110",
                      20 when "10101111111111",
                      20 when "10110000000000",
                      20 when "10110000000001",
                      20 when "10110000000010",
                      20 when "10110000000011",
                      20 when "10110000000100",
                      19 when "10110000000101",
                      19 when "10110000000110",
                      19 when "10110000000111",
                      19 when "10110000001000",
                      19 when "10110000001001",
                      19 when "10110000001010",
                      19 when "10110000001011",
                      19 when "10110000001100",
                      19 when "10110000001101",
                      19 when "10110000001110",
                      19 when "10110000001111",
                      19 when "10110000010000",
                      19 when "10110000010001",
                      19 when "10110000010010",
                      19 when "10110000010011",
                      19 when "10110000010100",
                      19 when "10110000010101",
                      19 when "10110000010110",
                      19 when "10110000010111",
                      19 when "10110000011000",
                      19 when "10110000011001",
                      19 when "10110000011010",
                      19 when "10110000011011",
                      19 when "10110000011100",
                      19 when "10110000011101",
                      19 when "10110000011110",
                      19 when "10110000011111",
                      19 when "10110000100000",
                      19 when "10110000100001",
                      19 when "10110000100010",
                      19 when "10110000100011",
                      19 when "10110000100100",
                      19 when "10110000100101",
                      19 when "10110000100110",
                      19 when "10110000100111",
                      19 when "10110000101000",
                      19 when "10110000101001",
                      19 when "10110000101010",
                      19 when "10110000101011",
                      19 when "10110000101100",
                      19 when "10110000101101",
                      19 when "10110000101110",
                      19 when "10110000101111",
                      19 when "10110000110000",
                      19 when "10110000110001",
                      19 when "10110000110010",
                      19 when "10110000110011",
                      19 when "10110000110100",
                      19 when "10110000110101",
                      19 when "10110000110110",
                      19 when "10110000110111",
                      19 when "10110000111000",
                      19 when "10110000111001",
                      19 when "10110000111010",
                      19 when "10110000111011",
                      19 when "10110000111100",
                      19 when "10110000111101",
                      19 when "10110000111110",
                      19 when "10110000111111",
                      19 when "10110001000000",
                      19 when "10110001000001",
                      19 when "10110001000010",
                      19 when "10110001000011",
                      19 when "10110001000100",
                      19 when "10110001000101",
                      19 when "10110001000110",
                      19 when "10110001000111",
                      19 when "10110001001000",
                      19 when "10110001001001",
                      19 when "10110001001010",
                      19 when "10110001001011",
                      19 when "10110001001100",
                      19 when "10110001001101",
                      19 when "10110001001110",
                      19 when "10110001001111",
                      19 when "10110001010000",
                      19 when "10110001010001",
                      19 when "10110001010010",
                      19 when "10110001010011",
                      19 when "10110001010100",
                      19 when "10110001010101",
                      19 when "10110001010110",
                      19 when "10110001010111",
                      19 when "10110001011000",
                      19 when "10110001011001",
                      19 when "10110001011010",
                      19 when "10110001011011",
                      19 when "10110001011100",
                      19 when "10110001011101",
                      19 when "10110001011110",
                      19 when "10110001011111",
                      19 when "10110001100000",
                      19 when "10110001100001",
                      19 when "10110001100010",
                      19 when "10110001100011",
                      19 when "10110001100100",
                      19 when "10110001100101",
                      19 when "10110001100110",
                      19 when "10110001100111",
                      19 when "10110001101000",
                      19 when "10110001101001",
                      19 when "10110001101010",
                      19 when "10110001101011",
                      19 when "10110001101100",
                      19 when "10110001101101",
                      19 when "10110001101110",
                      19 when "10110001101111",
                      19 when "10110001110000",
                      19 when "10110001110001",
                      19 when "10110001110010",
                      19 when "10110001110011",
                      19 when "10110001110100",
                      19 when "10110001110101",
                      19 when "10110001110110",
                      19 when "10110001110111",
                      19 when "10110001111000",
                      19 when "10110001111001",
                      19 when "10110001111010",
                      19 when "10110001111011",
                      19 when "10110001111100",
                      19 when "10110001111101",
                      19 when "10110001111110",
                      19 when "10110001111111",
                      19 when "10110010000000",
                      19 when "10110010000001",
                      19 when "10110010000010",
                      19 when "10110010000011",
                      19 when "10110010000100",
                      19 when "10110010000101",
                      19 when "10110010000110",
                      19 when "10110010000111",
                      19 when "10110010001000",
                      19 when "10110010001001",
                      19 when "10110010001010",
                      19 when "10110010001011",
                      19 when "10110010001100",
                      19 when "10110010001101",
                      19 when "10110010001110",
                      19 when "10110010001111",
                      19 when "10110010010000",
                      19 when "10110010010001",
                      19 when "10110010010010",
                      19 when "10110010010011",
                      19 when "10110010010100",
                      19 when "10110010010101",
                      19 when "10110010010110",
                      19 when "10110010010111",
                      19 when "10110010011000",
                      19 when "10110010011001",
                      19 when "10110010011010",
                      19 when "10110010011011",
                      19 when "10110010011100",
                      19 when "10110010011101",
                      19 when "10110010011110",
                      19 when "10110010011111",
                      19 when "10110010100000",
                      19 when "10110010100001",
                      19 when "10110010100010",
                      19 when "10110010100011",
                      19 when "10110010100100",
                      19 when "10110010100101",
                      19 when "10110010100110",
                      19 when "10110010100111",
                      19 when "10110010101000",
                      19 when "10110010101001",
                      19 when "10110010101010",
                      19 when "10110010101011",
                      19 when "10110010101100",
                      19 when "10110010101101",
                      19 when "10110010101110",
                      19 when "10110010101111",
                      19 when "10110010110000",
                      19 when "10110010110001",
                      19 when "10110010110010",
                      19 when "10110010110011",
                      19 when "10110010110100",
                      19 when "10110010110101",
                      19 when "10110010110110",
                      19 when "10110010110111",
                      19 when "10110010111000",
                      19 when "10110010111001",
                      19 when "10110010111010",
                      19 when "10110010111011",
                      19 when "10110010111100",
                      19 when "10110010111101",
                      19 when "10110010111110",
                      19 when "10110010111111",
                      19 when "10110011000000",
                      19 when "10110011000001",
                      19 when "10110011000010",
                      19 when "10110011000011",
                      19 when "10110011000100",
                      19 when "10110011000101",
                      19 when "10110011000110",
                      19 when "10110011000111",
                      19 when "10110011001000",
                      19 when "10110011001001",
                      19 when "10110011001010",
                      19 when "10110011001011",
                      19 when "10110011001100",
                      19 when "10110011001101",
                      19 when "10110011001110",
                      19 when "10110011001111",
                      19 when "10110011010000",
                      19 when "10110011010001",
                      19 when "10110011010010",
                      19 when "10110011010011",
                      19 when "10110011010100",
                      19 when "10110011010101",
                      19 when "10110011010110",
                      19 when "10110011010111",
                      19 when "10110011011000",
                      19 when "10110011011001",
                      19 when "10110011011010",
                      19 when "10110011011011",
                      19 when "10110011011100",
                      19 when "10110011011101",
                      19 when "10110011011110",
                      19 when "10110011011111",
                      19 when "10110011100000",
                      19 when "10110011100001",
                      19 when "10110011100010",
                      19 when "10110011100011",
                      19 when "10110011100100",
                      19 when "10110011100101",
                      19 when "10110011100110",
                      19 when "10110011100111",
                      19 when "10110011101000",
                      19 when "10110011101001",
                      19 when "10110011101010",
                      19 when "10110011101011",
                      19 when "10110011101100",
                      19 when "10110011101101",
                      19 when "10110011101110",
                      19 when "10110011101111",
                      19 when "10110011110000",
                      19 when "10110011110001",
                      19 when "10110011110010",
                      19 when "10110011110011",
                      19 when "10110011110100",
                      19 when "10110011110101",
                      19 when "10110011110110",
                      19 when "10110011110111",
                      19 when "10110011111000",
                      19 when "10110011111001",
                      19 when "10110011111010",
                      19 when "10110011111011",
                      19 when "10110011111100",
                      19 when "10110011111101",
                      19 when "10110011111110",
                      19 when "10110011111111",
                      19 when "10110100000000",
                      19 when "10110100000001",
                      19 when "10110100000010",
                      19 when "10110100000011",
                      19 when "10110100000100",
                      19 when "10110100000101",
                      19 when "10110100000110",
                      19 when "10110100000111",
                      19 when "10110100001000",
                      19 when "10110100001001",
                      19 when "10110100001010",
                      19 when "10110100001011",
                      19 when "10110100001100",
                      19 when "10110100001101",
                      19 when "10110100001110",
                      19 when "10110100001111",
                      19 when "10110100010000",
                      19 when "10110100010001",
                      19 when "10110100010010",
                      19 when "10110100010011",
                      19 when "10110100010100",
                      19 when "10110100010101",
                      19 when "10110100010110",
                      19 when "10110100010111",
                      19 when "10110100011000",
                      19 when "10110100011001",
                      19 when "10110100011010",
                      19 when "10110100011011",
                      19 when "10110100011100",
                      19 when "10110100011101",
                      19 when "10110100011110",
                      19 when "10110100011111",
                      19 when "10110100100000",
                      19 when "10110100100001",
                      19 when "10110100100010",
                      19 when "10110100100011",
                      19 when "10110100100100",
                      19 when "10110100100101",
                      19 when "10110100100110",
                      19 when "10110100100111",
                      19 when "10110100101000",
                      19 when "10110100101001",
                      19 when "10110100101010",
                      19 when "10110100101011",
                      19 when "10110100101100",
                      19 when "10110100101101",
                      19 when "10110100101110",
                      19 when "10110100101111",
                      19 when "10110100110000",
                      19 when "10110100110001",
                      19 when "10110100110010",
                      19 when "10110100110011",
                      19 when "10110100110100",
                      19 when "10110100110101",
                      19 when "10110100110110",
                      19 when "10110100110111",
                      19 when "10110100111000",
                      19 when "10110100111001",
                      19 when "10110100111010",
                      19 when "10110100111011",
                      19 when "10110100111100",
                      19 when "10110100111101",
                      19 when "10110100111110",
                      19 when "10110100111111",
                      19 when "10110101000000",
                      19 when "10110101000001",
                      19 when "10110101000010",
                      19 when "10110101000011",
                      19 when "10110101000100",
                      19 when "10110101000101",
                      19 when "10110101000110",
                      19 when "10110101000111",
                      19 when "10110101001000",
                      19 when "10110101001001",
                      19 when "10110101001010",
                      19 when "10110101001011",
                      19 when "10110101001100",
                      19 when "10110101001101",
                      19 when "10110101001110",
                      19 when "10110101001111",
                      19 when "10110101010000",
                      19 when "10110101010001",
                      19 when "10110101010010",
                      19 when "10110101010011",
                      19 when "10110101010100",
                      19 when "10110101010101",
                      19 when "10110101010110",
                      19 when "10110101010111",
                      19 when "10110101011000",
                      19 when "10110101011001",
                      19 when "10110101011010",
                      19 when "10110101011011",
                      19 when "10110101011100",
                      19 when "10110101011101",
                      19 when "10110101011110",
                      19 when "10110101011111",
                      19 when "10110101100000",
                      19 when "10110101100001",
                      19 when "10110101100010",
                      19 when "10110101100011",
                      19 when "10110101100100",
                      19 when "10110101100101",
                      19 when "10110101100110",
                      19 when "10110101100111",
                      19 when "10110101101000",
                      19 when "10110101101001",
                      19 when "10110101101010",
                      19 when "10110101101011",
                      19 when "10110101101100",
                      19 when "10110101101101",
                      19 when "10110101101110",
                      19 when "10110101101111",
                      19 when "10110101110000",
                      19 when "10110101110001",
                      19 when "10110101110010",
                      19 when "10110101110011",
                      19 when "10110101110100",
                      19 when "10110101110101",
                      19 when "10110101110110",
                      19 when "10110101110111",
                      19 when "10110101111000",
                      19 when "10110101111001",
                      19 when "10110101111010",
                      19 when "10110101111011",
                      19 when "10110101111100",
                      19 when "10110101111101",
                      19 when "10110101111110",
                      19 when "10110101111111",
                      19 when "10110110000000",
                      19 when "10110110000001",
                      19 when "10110110000010",
                      19 when "10110110000011",
                      19 when "10110110000100",
                      19 when "10110110000101",
                      19 when "10110110000110",
                      19 when "10110110000111",
                      19 when "10110110001000",
                      19 when "10110110001001",
                      19 when "10110110001010",
                      19 when "10110110001011",
                      19 when "10110110001100",
                      19 when "10110110001101",
                      19 when "10110110001110",
                      19 when "10110110001111",
                      19 when "10110110010000",
                      19 when "10110110010001",
                      19 when "10110110010010",
                      19 when "10110110010011",
                      19 when "10110110010100",
                      19 when "10110110010101",
                      19 when "10110110010110",
                      19 when "10110110010111",
                      19 when "10110110011000",
                      19 when "10110110011001",
                      19 when "10110110011010",
                      19 when "10110110011011",
                      19 when "10110110011100",
                      19 when "10110110011101",
                      19 when "10110110011110",
                      19 when "10110110011111",
                      19 when "10110110100000",
                      19 when "10110110100001",
                      19 when "10110110100010",
                      19 when "10110110100011",
                      19 when "10110110100100",
                      19 when "10110110100101",
                      19 when "10110110100110",
                      19 when "10110110100111",
                      19 when "10110110101000",
                      19 when "10110110101001",
                      19 when "10110110101010",
                      19 when "10110110101011",
                      19 when "10110110101100",
                      19 when "10110110101101",
                      19 when "10110110101110",
                      19 when "10110110101111",
                      19 when "10110110110000",
                      19 when "10110110110001",
                      19 when "10110110110010",
                      19 when "10110110110011",
                      19 when "10110110110100",
                      19 when "10110110110101",
                      19 when "10110110110110",
                      19 when "10110110110111",
                      19 when "10110110111000",
                      19 when "10110110111001",
                      19 when "10110110111010",
                      19 when "10110110111011",
                      19 when "10110110111100",
                      19 when "10110110111101",
                      19 when "10110110111110",
                      19 when "10110110111111",
                      19 when "10110111000000",
                      19 when "10110111000001",
                      19 when "10110111000010",
                      19 when "10110111000011",
                      19 when "10110111000100",
                      19 when "10110111000101",
                      19 when "10110111000110",
                      19 when "10110111000111",
                      19 when "10110111001000",
                      19 when "10110111001001",
                      19 when "10110111001010",
                      19 when "10110111001011",
                      19 when "10110111001100",
                      19 when "10110111001101",
                      19 when "10110111001110",
                      19 when "10110111001111",
                      19 when "10110111010000",
                      19 when "10110111010001",
                      19 when "10110111010010",
                      19 when "10110111010011",
                      19 when "10110111010100",
                      19 when "10110111010101",
                      19 when "10110111010110",
                      19 when "10110111010111",
                      19 when "10110111011000",
                      19 when "10110111011001",
                      19 when "10110111011010",
                      19 when "10110111011011",
                      19 when "10110111011100",
                      19 when "10110111011101",
                      19 when "10110111011110",
                      19 when "10110111011111",
                      19 when "10110111100000",
                      19 when "10110111100001",
                      19 when "10110111100010",
                      19 when "10110111100011",
                      19 when "10110111100100",
                      19 when "10110111100101",
                      19 when "10110111100110",
                      19 when "10110111100111",
                      19 when "10110111101000",
                      19 when "10110111101001",
                      19 when "10110111101010",
                      19 when "10110111101011",
                      19 when "10110111101100",
                      19 when "10110111101101",
                      19 when "10110111101110",
                      19 when "10110111101111",
                      19 when "10110111110000",
                      19 when "10110111110001",
                      19 when "10110111110010",
                      19 when "10110111110011",
                      19 when "10110111110100",
                      19 when "10110111110101",
                      19 when "10110111110110",
                      19 when "10110111110111",
                      19 when "10110111111000",
                      19 when "10110111111001",
                      19 when "10110111111010",
                      19 when "10110111111011",
                      19 when "10110111111100",
                      19 when "10110111111101",
                      19 when "10110111111110",
                      19 when "10110111111111",
                      19 when "10111000000000",
                      19 when "10111000000001",
                      19 when "10111000000010",
                      19 when "10111000000011",
                      19 when "10111000000100",
                      19 when "10111000000101",
                      19 when "10111000000110",
                      19 when "10111000000111",
                      19 when "10111000001000",
                      19 when "10111000001001",
                      19 when "10111000001010",
                      19 when "10111000001011",
                      19 when "10111000001100",
                      19 when "10111000001101",
                      19 when "10111000001110",
                      19 when "10111000001111",
                      19 when "10111000010000",
                      19 when "10111000010001",
                      19 when "10111000010010",
                      19 when "10111000010011",
                      19 when "10111000010100",
                      19 when "10111000010101",
                      19 when "10111000010110",
                      19 when "10111000010111",
                      19 when "10111000011000",
                      19 when "10111000011001",
                      19 when "10111000011010",
                      19 when "10111000011011",
                      19 when "10111000011100",
                      19 when "10111000011101",
                      19 when "10111000011110",
                      19 when "10111000011111",
                      19 when "10111000100000",
                      19 when "10111000100001",
                      19 when "10111000100010",
                      19 when "10111000100011",
                      19 when "10111000100100",
                      19 when "10111000100101",
                      19 when "10111000100110",
                      19 when "10111000100111",
                      19 when "10111000101000",
                      19 when "10111000101001",
                      19 when "10111000101010",
                      19 when "10111000101011",
                      19 when "10111000101100",
                      19 when "10111000101101",
                      19 when "10111000101110",
                      19 when "10111000101111",
                      19 when "10111000110000",
                      19 when "10111000110001",
                      19 when "10111000110010",
                      19 when "10111000110011",
                      19 when "10111000110100",
                      19 when "10111000110101",
                      19 when "10111000110110",
                      19 when "10111000110111",
                      19 when "10111000111000",
                      19 when "10111000111001",
                      19 when "10111000111010",
                      19 when "10111000111011",
                      19 when "10111000111100",
                      19 when "10111000111101",
                      19 when "10111000111110",
                      19 when "10111000111111",
                      19 when "10111001000000",
                      19 when "10111001000001",
                      19 when "10111001000010",
                      19 when "10111001000011",
                      19 when "10111001000100",
                      19 when "10111001000101",
                      19 when "10111001000110",
                      19 when "10111001000111",
                      19 when "10111001001000",
                      19 when "10111001001001",
                      19 when "10111001001010",
                      19 when "10111001001011",
                      19 when "10111001001100",
                      19 when "10111001001101",
                      19 when "10111001001110",
                      19 when "10111001001111",
                      19 when "10111001010000",
                      19 when "10111001010001",
                      19 when "10111001010010",
                      19 when "10111001010011",
                      19 when "10111001010100",
                      19 when "10111001010101",
                      19 when "10111001010110",
                      19 when "10111001010111",
                      19 when "10111001011000",
                      19 when "10111001011001",
                      19 when "10111001011010",
                      19 when "10111001011011",
                      19 when "10111001011100",
                      19 when "10111001011101",
                      19 when "10111001011110",
                      19 when "10111001011111",
                      19 when "10111001100000",
                      19 when "10111001100001",
                      19 when "10111001100010",
                      19 when "10111001100011",
                      19 when "10111001100100",
                      19 when "10111001100101",
                      18 when "10111001100110",
                      18 when "10111001100111",
                      18 when "10111001101000",
                      18 when "10111001101001",
                      18 when "10111001101010",
                      18 when "10111001101011",
                      18 when "10111001101100",
                      18 when "10111001101101",
                      18 when "10111001101110",
                      18 when "10111001101111",
                      18 when "10111001110000",
                      18 when "10111001110001",
                      18 when "10111001110010",
                      18 when "10111001110011",
                      18 when "10111001110100",
                      18 when "10111001110101",
                      18 when "10111001110110",
                      18 when "10111001110111",
                      18 when "10111001111000",
                      18 when "10111001111001",
                      18 when "10111001111010",
                      18 when "10111001111011",
                      18 when "10111001111100",
                      18 when "10111001111101",
                      18 when "10111001111110",
                      18 when "10111001111111",
                      18 when "10111010000000",
                      18 when "10111010000001",
                      18 when "10111010000010",
                      18 when "10111010000011",
                      18 when "10111010000100",
                      18 when "10111010000101",
                      18 when "10111010000110",
                      18 when "10111010000111",
                      18 when "10111010001000",
                      18 when "10111010001001",
                      18 when "10111010001010",
                      18 when "10111010001011",
                      18 when "10111010001100",
                      18 when "10111010001101",
                      18 when "10111010001110",
                      18 when "10111010001111",
                      18 when "10111010010000",
                      18 when "10111010010001",
                      18 when "10111010010010",
                      18 when "10111010010011",
                      18 when "10111010010100",
                      18 when "10111010010101",
                      18 when "10111010010110",
                      18 when "10111010010111",
                      18 when "10111010011000",
                      18 when "10111010011001",
                      18 when "10111010011010",
                      18 when "10111010011011",
                      18 when "10111010011100",
                      18 when "10111010011101",
                      18 when "10111010011110",
                      18 when "10111010011111",
                      18 when "10111010100000",
                      18 when "10111010100001",
                      18 when "10111010100010",
                      18 when "10111010100011",
                      18 when "10111010100100",
                      18 when "10111010100101",
                      18 when "10111010100110",
                      18 when "10111010100111",
                      18 when "10111010101000",
                      18 when "10111010101001",
                      18 when "10111010101010",
                      18 when "10111010101011",
                      18 when "10111010101100",
                      18 when "10111010101101",
                      18 when "10111010101110",
                      18 when "10111010101111",
                      18 when "10111010110000",
                      18 when "10111010110001",
                      18 when "10111010110010",
                      18 when "10111010110011",
                      18 when "10111010110100",
                      18 when "10111010110101",
                      18 when "10111010110110",
                      18 when "10111010110111",
                      18 when "10111010111000",
                      18 when "10111010111001",
                      18 when "10111010111010",
                      18 when "10111010111011",
                      18 when "10111010111100",
                      18 when "10111010111101",
                      18 when "10111010111110",
                      18 when "10111010111111",
                      18 when "10111011000000",
                      18 when "10111011000001",
                      18 when "10111011000010",
                      18 when "10111011000011",
                      18 when "10111011000100",
                      18 when "10111011000101",
                      18 when "10111011000110",
                      18 when "10111011000111",
                      18 when "10111011001000",
                      18 when "10111011001001",
                      18 when "10111011001010",
                      18 when "10111011001011",
                      18 when "10111011001100",
                      18 when "10111011001101",
                      18 when "10111011001110",
                      18 when "10111011001111",
                      18 when "10111011010000",
                      18 when "10111011010001",
                      18 when "10111011010010",
                      18 when "10111011010011",
                      18 when "10111011010100",
                      18 when "10111011010101",
                      18 when "10111011010110",
                      18 when "10111011010111",
                      18 when "10111011011000",
                      18 when "10111011011001",
                      18 when "10111011011010",
                      18 when "10111011011011",
                      18 when "10111011011100",
                      18 when "10111011011101",
                      18 when "10111011011110",
                      18 when "10111011011111",
                      18 when "10111011100000",
                      18 when "10111011100001",
                      18 when "10111011100010",
                      18 when "10111011100011",
                      18 when "10111011100100",
                      18 when "10111011100101",
                      18 when "10111011100110",
                      18 when "10111011100111",
                      18 when "10111011101000",
                      18 when "10111011101001",
                      18 when "10111011101010",
                      18 when "10111011101011",
                      18 when "10111011101100",
                      18 when "10111011101101",
                      18 when "10111011101110",
                      18 when "10111011101111",
                      18 when "10111011110000",
                      18 when "10111011110001",
                      18 when "10111011110010",
                      18 when "10111011110011",
                      18 when "10111011110100",
                      18 when "10111011110101",
                      18 when "10111011110110",
                      18 when "10111011110111",
                      18 when "10111011111000",
                      18 when "10111011111001",
                      18 when "10111011111010",
                      18 when "10111011111011",
                      18 when "10111011111100",
                      18 when "10111011111101",
                      18 when "10111011111110",
                      18 when "10111011111111",
                      18 when "10111100000000",
                      18 when "10111100000001",
                      18 when "10111100000010",
                      18 when "10111100000011",
                      18 when "10111100000100",
                      18 when "10111100000101",
                      18 when "10111100000110",
                      18 when "10111100000111",
                      18 when "10111100001000",
                      18 when "10111100001001",
                      18 when "10111100001010",
                      18 when "10111100001011",
                      18 when "10111100001100",
                      18 when "10111100001101",
                      18 when "10111100001110",
                      18 when "10111100001111",
                      18 when "10111100010000",
                      18 when "10111100010001",
                      18 when "10111100010010",
                      18 when "10111100010011",
                      18 when "10111100010100",
                      18 when "10111100010101",
                      18 when "10111100010110",
                      18 when "10111100010111",
                      18 when "10111100011000",
                      18 when "10111100011001",
                      18 when "10111100011010",
                      18 when "10111100011011",
                      18 when "10111100011100",
                      18 when "10111100011101",
                      18 when "10111100011110",
                      18 when "10111100011111",
                      18 when "10111100100000",
                      18 when "10111100100001",
                      18 when "10111100100010",
                      18 when "10111100100011",
                      18 when "10111100100100",
                      18 when "10111100100101",
                      18 when "10111100100110",
                      18 when "10111100100111",
                      18 when "10111100101000",
                      18 when "10111100101001",
                      18 when "10111100101010",
                      18 when "10111100101011",
                      18 when "10111100101100",
                      18 when "10111100101101",
                      18 when "10111100101110",
                      18 when "10111100101111",
                      18 when "10111100110000",
                      18 when "10111100110001",
                      18 when "10111100110010",
                      18 when "10111100110011",
                      18 when "10111100110100",
                      18 when "10111100110101",
                      18 when "10111100110110",
                      18 when "10111100110111",
                      18 when "10111100111000",
                      18 when "10111100111001",
                      18 when "10111100111010",
                      18 when "10111100111011",
                      18 when "10111100111100",
                      18 when "10111100111101",
                      18 when "10111100111110",
                      18 when "10111100111111",
                      18 when "10111101000000",
                      18 when "10111101000001",
                      18 when "10111101000010",
                      18 when "10111101000011",
                      18 when "10111101000100",
                      18 when "10111101000101",
                      18 when "10111101000110",
                      18 when "10111101000111",
                      18 when "10111101001000",
                      18 when "10111101001001",
                      18 when "10111101001010",
                      18 when "10111101001011",
                      18 when "10111101001100",
                      18 when "10111101001101",
                      18 when "10111101001110",
                      18 when "10111101001111",
                      18 when "10111101010000",
                      18 when "10111101010001",
                      18 when "10111101010010",
                      18 when "10111101010011",
                      18 when "10111101010100",
                      18 when "10111101010101",
                      18 when "10111101010110",
                      18 when "10111101010111",
                      18 when "10111101011000",
                      18 when "10111101011001",
                      18 when "10111101011010",
                      18 when "10111101011011",
                      18 when "10111101011100",
                      18 when "10111101011101",
                      18 when "10111101011110",
                      18 when "10111101011111",
                      18 when "10111101100000",
                      18 when "10111101100001",
                      18 when "10111101100010",
                      18 when "10111101100011",
                      18 when "10111101100100",
                      18 when "10111101100101",
                      18 when "10111101100110",
                      18 when "10111101100111",
                      18 when "10111101101000",
                      18 when "10111101101001",
                      18 when "10111101101010",
                      18 when "10111101101011",
                      18 when "10111101101100",
                      18 when "10111101101101",
                      18 when "10111101101110",
                      18 when "10111101101111",
                      18 when "10111101110000",
                      18 when "10111101110001",
                      18 when "10111101110010",
                      18 when "10111101110011",
                      18 when "10111101110100",
                      18 when "10111101110101",
                      18 when "10111101110110",
                      18 when "10111101110111",
                      18 when "10111101111000",
                      18 when "10111101111001",
                      18 when "10111101111010",
                      18 when "10111101111011",
                      18 when "10111101111100",
                      18 when "10111101111101",
                      18 when "10111101111110",
                      18 when "10111101111111",
                      18 when "10111110000000",
                      18 when "10111110000001",
                      18 when "10111110000010",
                      18 when "10111110000011",
                      18 when "10111110000100",
                      18 when "10111110000101",
                      18 when "10111110000110",
                      18 when "10111110000111",
                      18 when "10111110001000",
                      18 when "10111110001001",
                      18 when "10111110001010",
                      18 when "10111110001011",
                      18 when "10111110001100",
                      18 when "10111110001101",
                      18 when "10111110001110",
                      18 when "10111110001111",
                      18 when "10111110010000",
                      18 when "10111110010001",
                      18 when "10111110010010",
                      18 when "10111110010011",
                      18 when "10111110010100",
                      18 when "10111110010101",
                      18 when "10111110010110",
                      18 when "10111110010111",
                      18 when "10111110011000",
                      18 when "10111110011001",
                      18 when "10111110011010",
                      18 when "10111110011011",
                      18 when "10111110011100",
                      18 when "10111110011101",
                      18 when "10111110011110",
                      18 when "10111110011111",
                      18 when "10111110100000",
                      18 when "10111110100001",
                      18 when "10111110100010",
                      18 when "10111110100011",
                      18 when "10111110100100",
                      18 when "10111110100101",
                      18 when "10111110100110",
                      18 when "10111110100111",
                      18 when "10111110101000",
                      18 when "10111110101001",
                      18 when "10111110101010",
                      18 when "10111110101011",
                      18 when "10111110101100",
                      18 when "10111110101101",
                      18 when "10111110101110",
                      18 when "10111110101111",
                      18 when "10111110110000",
                      18 when "10111110110001",
                      18 when "10111110110010",
                      18 when "10111110110011",
                      18 when "10111110110100",
                      18 when "10111110110101",
                      18 when "10111110110110",
                      18 when "10111110110111",
                      18 when "10111110111000",
                      18 when "10111110111001",
                      18 when "10111110111010",
                      18 when "10111110111011",
                      18 when "10111110111100",
                      18 when "10111110111101",
                      18 when "10111110111110",
                      18 when "10111110111111",
                      18 when "10111111000000",
                      18 when "10111111000001",
                      18 when "10111111000010",
                      18 when "10111111000011",
                      18 when "10111111000100",
                      18 when "10111111000101",
                      18 when "10111111000110",
                      18 when "10111111000111",
                      18 when "10111111001000",
                      18 when "10111111001001",
                      18 when "10111111001010",
                      18 when "10111111001011",
                      18 when "10111111001100",
                      18 when "10111111001101",
                      18 when "10111111001110",
                      18 when "10111111001111",
                      18 when "10111111010000",
                      18 when "10111111010001",
                      18 when "10111111010010",
                      18 when "10111111010011",
                      18 when "10111111010100",
                      18 when "10111111010101",
                      18 when "10111111010110",
                      18 when "10111111010111",
                      18 when "10111111011000",
                      18 when "10111111011001",
                      18 when "10111111011010",
                      18 when "10111111011011",
                      18 when "10111111011100",
                      18 when "10111111011101",
                      18 when "10111111011110",
                      18 when "10111111011111",
                      18 when "10111111100000",
                      18 when "10111111100001",
                      18 when "10111111100010",
                      18 when "10111111100011",
                      18 when "10111111100100",
                      18 when "10111111100101",
                      18 when "10111111100110",
                      18 when "10111111100111",
                      18 when "10111111101000",
                      18 when "10111111101001",
                      18 when "10111111101010",
                      18 when "10111111101011",
                      18 when "10111111101100",
                      18 when "10111111101101",
                      18 when "10111111101110",
                      18 when "10111111101111",
                      18 when "10111111110000",
                      18 when "10111111110001",
                      18 when "10111111110010",
                      18 when "10111111110011",
                      18 when "10111111110100",
                      18 when "10111111110101",
                      18 when "10111111110110",
                      18 when "10111111110111",
                      18 when "10111111111000",
                      18 when "10111111111001",
                      18 when "10111111111010",
                      18 when "10111111111011",
                      18 when "10111111111100",
                      18 when "10111111111101",
                      18 when "10111111111110",
                      18 when "10111111111111",
                      18 when "11000000000000",
                      18 when "11000000000001",
                      18 when "11000000000010",
                      18 when "11000000000011",
                      18 when "11000000000100",
                      18 when "11000000000101",
                      18 when "11000000000110",
                      18 when "11000000000111",
                      18 when "11000000001000",
                      18 when "11000000001001",
                      18 when "11000000001010",
                      18 when "11000000001011",
                      18 when "11000000001100",
                      18 when "11000000001101",
                      18 when "11000000001110",
                      18 when "11000000001111",
                      18 when "11000000010000",
                      18 when "11000000010001",
                      18 when "11000000010010",
                      18 when "11000000010011",
                      18 when "11000000010100",
                      18 when "11000000010101",
                      18 when "11000000010110",
                      18 when "11000000010111",
                      18 when "11000000011000",
                      18 when "11000000011001",
                      18 when "11000000011010",
                      18 when "11000000011011",
                      18 when "11000000011100",
                      18 when "11000000011101",
                      18 when "11000000011110",
                      18 when "11000000011111",
                      18 when "11000000100000",
                      18 when "11000000100001",
                      18 when "11000000100010",
                      18 when "11000000100011",
                      18 when "11000000100100",
                      18 when "11000000100101",
                      18 when "11000000100110",
                      18 when "11000000100111",
                      18 when "11000000101000",
                      18 when "11000000101001",
                      18 when "11000000101010",
                      18 when "11000000101011",
                      18 when "11000000101100",
                      18 when "11000000101101",
                      18 when "11000000101110",
                      18 when "11000000101111",
                      18 when "11000000110000",
                      18 when "11000000110001",
                      18 when "11000000110010",
                      18 when "11000000110011",
                      18 when "11000000110100",
                      18 when "11000000110101",
                      18 when "11000000110110",
                      18 when "11000000110111",
                      18 when "11000000111000",
                      18 when "11000000111001",
                      18 when "11000000111010",
                      18 when "11000000111011",
                      18 when "11000000111100",
                      18 when "11000000111101",
                      18 when "11000000111110",
                      18 when "11000000111111",
                      18 when "11000001000000",
                      18 when "11000001000001",
                      18 when "11000001000010",
                      18 when "11000001000011",
                      18 when "11000001000100",
                      18 when "11000001000101",
                      18 when "11000001000110",
                      18 when "11000001000111",
                      18 when "11000001001000",
                      18 when "11000001001001",
                      18 when "11000001001010",
                      18 when "11000001001011",
                      18 when "11000001001100",
                      18 when "11000001001101",
                      18 when "11000001001110",
                      18 when "11000001001111",
                      18 when "11000001010000",
                      18 when "11000001010001",
                      18 when "11000001010010",
                      18 when "11000001010011",
                      18 when "11000001010100",
                      18 when "11000001010101",
                      18 when "11000001010110",
                      18 when "11000001010111",
                      18 when "11000001011000",
                      18 when "11000001011001",
                      18 when "11000001011010",
                      18 when "11000001011011",
                      18 when "11000001011100",
                      18 when "11000001011101",
                      18 when "11000001011110",
                      18 when "11000001011111",
                      18 when "11000001100000",
                      18 when "11000001100001",
                      18 when "11000001100010",
                      18 when "11000001100011",
                      18 when "11000001100100",
                      18 when "11000001100101",
                      18 when "11000001100110",
                      18 when "11000001100111",
                      18 when "11000001101000",
                      18 when "11000001101001",
                      18 when "11000001101010",
                      18 when "11000001101011",
                      18 when "11000001101100",
                      18 when "11000001101101",
                      18 when "11000001101110",
                      18 when "11000001101111",
                      18 when "11000001110000",
                      18 when "11000001110001",
                      18 when "11000001110010",
                      18 when "11000001110011",
                      18 when "11000001110100",
                      18 when "11000001110101",
                      18 when "11000001110110",
                      18 when "11000001110111",
                      18 when "11000001111000",
                      18 when "11000001111001",
                      18 when "11000001111010",
                      18 when "11000001111011",
                      18 when "11000001111100",
                      18 when "11000001111101",
                      18 when "11000001111110",
                      18 when "11000001111111",
                      18 when "11000010000000",
                      18 when "11000010000001",
                      18 when "11000010000010",
                      18 when "11000010000011",
                      18 when "11000010000100",
                      18 when "11000010000101",
                      18 when "11000010000110",
                      18 when "11000010000111",
                      18 when "11000010001000",
                      18 when "11000010001001",
                      18 when "11000010001010",
                      18 when "11000010001011",
                      18 when "11000010001100",
                      18 when "11000010001101",
                      18 when "11000010001110",
                      18 when "11000010001111",
                      18 when "11000010010000",
                      18 when "11000010010001",
                      18 when "11000010010010",
                      18 when "11000010010011",
                      18 when "11000010010100",
                      18 when "11000010010101",
                      18 when "11000010010110",
                      18 when "11000010010111",
                      18 when "11000010011000",
                      18 when "11000010011001",
                      18 when "11000010011010",
                      18 when "11000010011011",
                      18 when "11000010011100",
                      18 when "11000010011101",
                      18 when "11000010011110",
                      18 when "11000010011111",
                      18 when "11000010100000",
                      18 when "11000010100001",
                      18 when "11000010100010",
                      18 when "11000010100011",
                      18 when "11000010100100",
                      18 when "11000010100101",
                      18 when "11000010100110",
                      18 when "11000010100111",
                      18 when "11000010101000",
                      18 when "11000010101001",
                      18 when "11000010101010",
                      18 when "11000010101011",
                      18 when "11000010101100",
                      18 when "11000010101101",
                      18 when "11000010101110",
                      18 when "11000010101111",
                      18 when "11000010110000",
                      18 when "11000010110001",
                      18 when "11000010110010",
                      18 when "11000010110011",
                      18 when "11000010110100",
                      18 when "11000010110101",
                      18 when "11000010110110",
                      18 when "11000010110111",
                      18 when "11000010111000",
                      18 when "11000010111001",
                      18 when "11000010111010",
                      18 when "11000010111011",
                      18 when "11000010111100",
                      18 when "11000010111101",
                      18 when "11000010111110",
                      18 when "11000010111111",
                      18 when "11000011000000",
                      18 when "11000011000001",
                      18 when "11000011000010",
                      18 when "11000011000011",
                      18 when "11000011000100",
                      18 when "11000011000101",
                      18 when "11000011000110",
                      18 when "11000011000111",
                      18 when "11000011001000",
                      18 when "11000011001001",
                      18 when "11000011001010",
                      18 when "11000011001011",
                      18 when "11000011001100",
                      18 when "11000011001101",
                      18 when "11000011001110",
                      18 when "11000011001111",
                      18 when "11000011010000",
                      18 when "11000011010001",
                      18 when "11000011010010",
                      18 when "11000011010011",
                      18 when "11000011010100",
                      18 when "11000011010101",
                      18 when "11000011010110",
                      18 when "11000011010111",
                      18 when "11000011011000",
                      18 when "11000011011001",
                      18 when "11000011011010",
                      18 when "11000011011011",
                      18 when "11000011011100",
                      18 when "11000011011101",
                      18 when "11000011011110",
                      18 when "11000011011111",
                      18 when "11000011100000",
                      18 when "11000011100001",
                      18 when "11000011100010",
                      18 when "11000011100011",
                      18 when "11000011100100",
                      18 when "11000011100101",
                      18 when "11000011100110",
                      18 when "11000011100111",
                      18 when "11000011101000",
                      18 when "11000011101001",
                      18 when "11000011101010",
                      18 when "11000011101011",
                      18 when "11000011101100",
                      18 when "11000011101101",
                      18 when "11000011101110",
                      18 when "11000011101111",
                      18 when "11000011110000",
                      18 when "11000011110001",
                      18 when "11000011110010",
                      18 when "11000011110011",
                      18 when "11000011110100",
                      18 when "11000011110101",
                      18 when "11000011110110",
                      18 when "11000011110111",
                      18 when "11000011111000",
                      18 when "11000011111001",
                      18 when "11000011111010",
                      18 when "11000011111011",
                      18 when "11000011111100",
                      18 when "11000011111101",
                      18 when "11000011111110",
                      18 when "11000011111111",
                      18 when "11000100000000",
                      18 when "11000100000001",
                      18 when "11000100000010",
                      18 when "11000100000011",
                      18 when "11000100000100",
                      18 when "11000100000101",
                      18 when "11000100000110",
                      18 when "11000100000111",
                      18 when "11000100001000",
                      18 when "11000100001001",
                      18 when "11000100001010",
                      18 when "11000100001011",
                      17 when "11000100001100",
                      17 when "11000100001101",
                      17 when "11000100001110",
                      17 when "11000100001111",
                      17 when "11000100010000",
                      17 when "11000100010001",
                      17 when "11000100010010",
                      17 when "11000100010011",
                      17 when "11000100010100",
                      17 when "11000100010101",
                      17 when "11000100010110",
                      17 when "11000100010111",
                      17 when "11000100011000",
                      17 when "11000100011001",
                      17 when "11000100011010",
                      17 when "11000100011011",
                      17 when "11000100011100",
                      17 when "11000100011101",
                      17 when "11000100011110",
                      17 when "11000100011111",
                      17 when "11000100100000",
                      17 when "11000100100001",
                      17 when "11000100100010",
                      17 when "11000100100011",
                      17 when "11000100100100",
                      17 when "11000100100101",
                      17 when "11000100100110",
                      17 when "11000100100111",
                      17 when "11000100101000",
                      17 when "11000100101001",
                      17 when "11000100101010",
                      17 when "11000100101011",
                      17 when "11000100101100",
                      17 when "11000100101101",
                      17 when "11000100101110",
                      17 when "11000100101111",
                      17 when "11000100110000",
                      17 when "11000100110001",
                      17 when "11000100110010",
                      17 when "11000100110011",
                      17 when "11000100110100",
                      17 when "11000100110101",
                      17 when "11000100110110",
                      17 when "11000100110111",
                      17 when "11000100111000",
                      17 when "11000100111001",
                      17 when "11000100111010",
                      17 when "11000100111011",
                      17 when "11000100111100",
                      17 when "11000100111101",
                      17 when "11000100111110",
                      17 when "11000100111111",
                      17 when "11000101000000",
                      17 when "11000101000001",
                      17 when "11000101000010",
                      17 when "11000101000011",
                      17 when "11000101000100",
                      17 when "11000101000101",
                      17 when "11000101000110",
                      17 when "11000101000111",
                      17 when "11000101001000",
                      17 when "11000101001001",
                      17 when "11000101001010",
                      17 when "11000101001011",
                      17 when "11000101001100",
                      17 when "11000101001101",
                      17 when "11000101001110",
                      17 when "11000101001111",
                      17 when "11000101010000",
                      17 when "11000101010001",
                      17 when "11000101010010",
                      17 when "11000101010011",
                      17 when "11000101010100",
                      17 when "11000101010101",
                      17 when "11000101010110",
                      17 when "11000101010111",
                      17 when "11000101011000",
                      17 when "11000101011001",
                      17 when "11000101011010",
                      17 when "11000101011011",
                      17 when "11000101011100",
                      17 when "11000101011101",
                      17 when "11000101011110",
                      17 when "11000101011111",
                      17 when "11000101100000",
                      17 when "11000101100001",
                      17 when "11000101100010",
                      17 when "11000101100011",
                      17 when "11000101100100",
                      17 when "11000101100101",
                      17 when "11000101100110",
                      17 when "11000101100111",
                      17 when "11000101101000",
                      17 when "11000101101001",
                      17 when "11000101101010",
                      17 when "11000101101011",
                      17 when "11000101101100",
                      17 when "11000101101101",
                      17 when "11000101101110",
                      17 when "11000101101111",
                      17 when "11000101110000",
                      17 when "11000101110001",
                      17 when "11000101110010",
                      17 when "11000101110011",
                      17 when "11000101110100",
                      17 when "11000101110101",
                      17 when "11000101110110",
                      17 when "11000101110111",
                      17 when "11000101111000",
                      17 when "11000101111001",
                      17 when "11000101111010",
                      17 when "11000101111011",
                      17 when "11000101111100",
                      17 when "11000101111101",
                      17 when "11000101111110",
                      17 when "11000101111111",
                      17 when "11000110000000",
                      17 when "11000110000001",
                      17 when "11000110000010",
                      17 when "11000110000011",
                      17 when "11000110000100",
                      17 when "11000110000101",
                      17 when "11000110000110",
                      17 when "11000110000111",
                      17 when "11000110001000",
                      17 when "11000110001001",
                      17 when "11000110001010",
                      17 when "11000110001011",
                      17 when "11000110001100",
                      17 when "11000110001101",
                      17 when "11000110001110",
                      17 when "11000110001111",
                      17 when "11000110010000",
                      17 when "11000110010001",
                      17 when "11000110010010",
                      17 when "11000110010011",
                      17 when "11000110010100",
                      17 when "11000110010101",
                      17 when "11000110010110",
                      17 when "11000110010111",
                      17 when "11000110011000",
                      17 when "11000110011001",
                      17 when "11000110011010",
                      17 when "11000110011011",
                      17 when "11000110011100",
                      17 when "11000110011101",
                      17 when "11000110011110",
                      17 when "11000110011111",
                      17 when "11000110100000",
                      17 when "11000110100001",
                      17 when "11000110100010",
                      17 when "11000110100011",
                      17 when "11000110100100",
                      17 when "11000110100101",
                      17 when "11000110100110",
                      17 when "11000110100111",
                      17 when "11000110101000",
                      17 when "11000110101001",
                      17 when "11000110101010",
                      17 when "11000110101011",
                      17 when "11000110101100",
                      17 when "11000110101101",
                      17 when "11000110101110",
                      17 when "11000110101111",
                      17 when "11000110110000",
                      17 when "11000110110001",
                      17 when "11000110110010",
                      17 when "11000110110011",
                      17 when "11000110110100",
                      17 when "11000110110101",
                      17 when "11000110110110",
                      17 when "11000110110111",
                      17 when "11000110111000",
                      17 when "11000110111001",
                      17 when "11000110111010",
                      17 when "11000110111011",
                      17 when "11000110111100",
                      17 when "11000110111101",
                      17 when "11000110111110",
                      17 when "11000110111111",
                      17 when "11000111000000",
                      17 when "11000111000001",
                      17 when "11000111000010",
                      17 when "11000111000011",
                      17 when "11000111000100",
                      17 when "11000111000101",
                      17 when "11000111000110",
                      17 when "11000111000111",
                      17 when "11000111001000",
                      17 when "11000111001001",
                      17 when "11000111001010",
                      17 when "11000111001011",
                      17 when "11000111001100",
                      17 when "11000111001101",
                      17 when "11000111001110",
                      17 when "11000111001111",
                      17 when "11000111010000",
                      17 when "11000111010001",
                      17 when "11000111010010",
                      17 when "11000111010011",
                      17 when "11000111010100",
                      17 when "11000111010101",
                      17 when "11000111010110",
                      17 when "11000111010111",
                      17 when "11000111011000",
                      17 when "11000111011001",
                      17 when "11000111011010",
                      17 when "11000111011011",
                      17 when "11000111011100",
                      17 when "11000111011101",
                      17 when "11000111011110",
                      17 when "11000111011111",
                      17 when "11000111100000",
                      17 when "11000111100001",
                      17 when "11000111100010",
                      17 when "11000111100011",
                      17 when "11000111100100",
                      17 when "11000111100101",
                      17 when "11000111100110",
                      17 when "11000111100111",
                      17 when "11000111101000",
                      17 when "11000111101001",
                      17 when "11000111101010",
                      17 when "11000111101011",
                      17 when "11000111101100",
                      17 when "11000111101101",
                      17 when "11000111101110",
                      17 when "11000111101111",
                      17 when "11000111110000",
                      17 when "11000111110001",
                      17 when "11000111110010",
                      17 when "11000111110011",
                      17 when "11000111110100",
                      17 when "11000111110101",
                      17 when "11000111110110",
                      17 when "11000111110111",
                      17 when "11000111111000",
                      17 when "11000111111001",
                      17 when "11000111111010",
                      17 when "11000111111011",
                      17 when "11000111111100",
                      17 when "11000111111101",
                      17 when "11000111111110",
                      17 when "11000111111111",
                      17 when "11001000000000",
                      17 when "11001000000001",
                      17 when "11001000000010",
                      17 when "11001000000011",
                      17 when "11001000000100",
                      17 when "11001000000101",
                      17 when "11001000000110",
                      17 when "11001000000111",
                      17 when "11001000001000",
                      17 when "11001000001001",
                      17 when "11001000001010",
                      17 when "11001000001011",
                      17 when "11001000001100",
                      17 when "11001000001101",
                      17 when "11001000001110",
                      17 when "11001000001111",
                      17 when "11001000010000",
                      17 when "11001000010001",
                      17 when "11001000010010",
                      17 when "11001000010011",
                      17 when "11001000010100",
                      17 when "11001000010101",
                      17 when "11001000010110",
                      17 when "11001000010111",
                      17 when "11001000011000",
                      17 when "11001000011001",
                      17 when "11001000011010",
                      17 when "11001000011011",
                      17 when "11001000011100",
                      17 when "11001000011101",
                      17 when "11001000011110",
                      17 when "11001000011111",
                      17 when "11001000100000",
                      17 when "11001000100001",
                      17 when "11001000100010",
                      17 when "11001000100011",
                      17 when "11001000100100",
                      17 when "11001000100101",
                      17 when "11001000100110",
                      17 when "11001000100111",
                      17 when "11001000101000",
                      17 when "11001000101001",
                      17 when "11001000101010",
                      17 when "11001000101011",
                      17 when "11001000101100",
                      17 when "11001000101101",
                      17 when "11001000101110",
                      17 when "11001000101111",
                      17 when "11001000110000",
                      17 when "11001000110001",
                      17 when "11001000110010",
                      17 when "11001000110011",
                      17 when "11001000110100",
                      17 when "11001000110101",
                      17 when "11001000110110",
                      17 when "11001000110111",
                      17 when "11001000111000",
                      17 when "11001000111001",
                      17 when "11001000111010",
                      17 when "11001000111011",
                      17 when "11001000111100",
                      17 when "11001000111101",
                      17 when "11001000111110",
                      17 when "11001000111111",
                      17 when "11001001000000",
                      17 when "11001001000001",
                      17 when "11001001000010",
                      17 when "11001001000011",
                      17 when "11001001000100",
                      17 when "11001001000101",
                      17 when "11001001000110",
                      17 when "11001001000111",
                      17 when "11001001001000",
                      17 when "11001001001001",
                      17 when "11001001001010",
                      17 when "11001001001011",
                      17 when "11001001001100",
                      17 when "11001001001101",
                      17 when "11001001001110",
                      17 when "11001001001111",
                      17 when "11001001010000",
                      17 when "11001001010001",
                      17 when "11001001010010",
                      17 when "11001001010011",
                      17 when "11001001010100",
                      17 when "11001001010101",
                      17 when "11001001010110",
                      17 when "11001001010111",
                      17 when "11001001011000",
                      17 when "11001001011001",
                      17 when "11001001011010",
                      17 when "11001001011011",
                      17 when "11001001011100",
                      17 when "11001001011101",
                      17 when "11001001011110",
                      17 when "11001001011111",
                      17 when "11001001100000",
                      17 when "11001001100001",
                      17 when "11001001100010",
                      17 when "11001001100011",
                      17 when "11001001100100",
                      17 when "11001001100101",
                      17 when "11001001100110",
                      17 when "11001001100111",
                      17 when "11001001101000",
                      17 when "11001001101001",
                      17 when "11001001101010",
                      17 when "11001001101011",
                      17 when "11001001101100",
                      17 when "11001001101101",
                      17 when "11001001101110",
                      17 when "11001001101111",
                      17 when "11001001110000",
                      17 when "11001001110001",
                      17 when "11001001110010",
                      17 when "11001001110011",
                      17 when "11001001110100",
                      17 when "11001001110101",
                      17 when "11001001110110",
                      17 when "11001001110111",
                      17 when "11001001111000",
                      17 when "11001001111001",
                      17 when "11001001111010",
                      17 when "11001001111011",
                      17 when "11001001111100",
                      17 when "11001001111101",
                      17 when "11001001111110",
                      17 when "11001001111111",
                      17 when "11001010000000",
                      17 when "11001010000001",
                      17 when "11001010000010",
                      17 when "11001010000011",
                      17 when "11001010000100",
                      17 when "11001010000101",
                      17 when "11001010000110",
                      17 when "11001010000111",
                      17 when "11001010001000",
                      17 when "11001010001001",
                      17 when "11001010001010",
                      17 when "11001010001011",
                      17 when "11001010001100",
                      17 when "11001010001101",
                      17 when "11001010001110",
                      17 when "11001010001111",
                      17 when "11001010010000",
                      17 when "11001010010001",
                      17 when "11001010010010",
                      17 when "11001010010011",
                      17 when "11001010010100",
                      17 when "11001010010101",
                      17 when "11001010010110",
                      17 when "11001010010111",
                      17 when "11001010011000",
                      17 when "11001010011001",
                      17 when "11001010011010",
                      17 when "11001010011011",
                      17 when "11001010011100",
                      17 when "11001010011101",
                      17 when "11001010011110",
                      17 when "11001010011111",
                      17 when "11001010100000",
                      17 when "11001010100001",
                      17 when "11001010100010",
                      17 when "11001010100011",
                      17 when "11001010100100",
                      17 when "11001010100101",
                      17 when "11001010100110",
                      17 when "11001010100111",
                      17 when "11001010101000",
                      17 when "11001010101001",
                      17 when "11001010101010",
                      17 when "11001010101011",
                      17 when "11001010101100",
                      17 when "11001010101101",
                      17 when "11001010101110",
                      17 when "11001010101111",
                      17 when "11001010110000",
                      17 when "11001010110001",
                      17 when "11001010110010",
                      17 when "11001010110011",
                      17 when "11001010110100",
                      17 when "11001010110101",
                      17 when "11001010110110",
                      17 when "11001010110111",
                      17 when "11001010111000",
                      17 when "11001010111001",
                      17 when "11001010111010",
                      17 when "11001010111011",
                      17 when "11001010111100",
                      17 when "11001010111101",
                      17 when "11001010111110",
                      17 when "11001010111111",
                      17 when "11001011000000",
                      17 when "11001011000001",
                      17 when "11001011000010",
                      17 when "11001011000011",
                      17 when "11001011000100",
                      17 when "11001011000101",
                      17 when "11001011000110",
                      17 when "11001011000111",
                      17 when "11001011001000",
                      17 when "11001011001001",
                      17 when "11001011001010",
                      17 when "11001011001011",
                      17 when "11001011001100",
                      17 when "11001011001101",
                      17 when "11001011001110",
                      17 when "11001011001111",
                      17 when "11001011010000",
                      17 when "11001011010001",
                      17 when "11001011010010",
                      17 when "11001011010011",
                      17 when "11001011010100",
                      17 when "11001011010101",
                      17 when "11001011010110",
                      17 when "11001011010111",
                      17 when "11001011011000",
                      17 when "11001011011001",
                      17 when "11001011011010",
                      17 when "11001011011011",
                      17 when "11001011011100",
                      17 when "11001011011101",
                      17 when "11001011011110",
                      17 when "11001011011111",
                      17 when "11001011100000",
                      17 when "11001011100001",
                      17 when "11001011100010",
                      17 when "11001011100011",
                      17 when "11001011100100",
                      17 when "11001011100101",
                      17 when "11001011100110",
                      17 when "11001011100111",
                      17 when "11001011101000",
                      17 when "11001011101001",
                      17 when "11001011101010",
                      17 when "11001011101011",
                      17 when "11001011101100",
                      17 when "11001011101101",
                      17 when "11001011101110",
                      17 when "11001011101111",
                      17 when "11001011110000",
                      17 when "11001011110001",
                      17 when "11001011110010",
                      17 when "11001011110011",
                      17 when "11001011110100",
                      17 when "11001011110101",
                      17 when "11001011110110",
                      17 when "11001011110111",
                      17 when "11001011111000",
                      17 when "11001011111001",
                      17 when "11001011111010",
                      17 when "11001011111011",
                      17 when "11001011111100",
                      17 when "11001011111101",
                      17 when "11001011111110",
                      17 when "11001011111111",
                      17 when "11001100000000",
                      17 when "11001100000001",
                      17 when "11001100000010",
                      17 when "11001100000011",
                      17 when "11001100000100",
                      17 when "11001100000101",
                      17 when "11001100000110",
                      17 when "11001100000111",
                      17 when "11001100001000",
                      17 when "11001100001001",
                      17 when "11001100001010",
                      17 when "11001100001011",
                      17 when "11001100001100",
                      17 when "11001100001101",
                      17 when "11001100001110",
                      17 when "11001100001111",
                      17 when "11001100010000",
                      17 when "11001100010001",
                      17 when "11001100010010",
                      17 when "11001100010011",
                      17 when "11001100010100",
                      17 when "11001100010101",
                      17 when "11001100010110",
                      17 when "11001100010111",
                      17 when "11001100011000",
                      17 when "11001100011001",
                      17 when "11001100011010",
                      17 when "11001100011011",
                      17 when "11001100011100",
                      17 when "11001100011101",
                      17 when "11001100011110",
                      17 when "11001100011111",
                      17 when "11001100100000",
                      17 when "11001100100001",
                      17 when "11001100100010",
                      17 when "11001100100011",
                      17 when "11001100100100",
                      17 when "11001100100101",
                      17 when "11001100100110",
                      17 when "11001100100111",
                      17 when "11001100101000",
                      17 when "11001100101001",
                      17 when "11001100101010",
                      17 when "11001100101011",
                      17 when "11001100101100",
                      17 when "11001100101101",
                      17 when "11001100101110",
                      17 when "11001100101111",
                      17 when "11001100110000",
                      17 when "11001100110001",
                      17 when "11001100110010",
                      17 when "11001100110011",
                      17 when "11001100110100",
                      17 when "11001100110101",
                      17 when "11001100110110",
                      17 when "11001100110111",
                      17 when "11001100111000",
                      17 when "11001100111001",
                      17 when "11001100111010",
                      17 when "11001100111011",
                      17 when "11001100111100",
                      17 when "11001100111101",
                      17 when "11001100111110",
                      17 when "11001100111111",
                      17 when "11001101000000",
                      17 when "11001101000001",
                      17 when "11001101000010",
                      17 when "11001101000011",
                      17 when "11001101000100",
                      17 when "11001101000101",
                      17 when "11001101000110",
                      17 when "11001101000111",
                      17 when "11001101001000",
                      17 when "11001101001001",
                      17 when "11001101001010",
                      17 when "11001101001011",
                      17 when "11001101001100",
                      17 when "11001101001101",
                      17 when "11001101001110",
                      17 when "11001101001111",
                      17 when "11001101010000",
                      17 when "11001101010001",
                      17 when "11001101010010",
                      17 when "11001101010011",
                      17 when "11001101010100",
                      17 when "11001101010101",
                      17 when "11001101010110",
                      17 when "11001101010111",
                      17 when "11001101011000",
                      17 when "11001101011001",
                      17 when "11001101011010",
                      17 when "11001101011011",
                      17 when "11001101011100",
                      17 when "11001101011101",
                      17 when "11001101011110",
                      17 when "11001101011111",
                      17 when "11001101100000",
                      17 when "11001101100001",
                      17 when "11001101100010",
                      17 when "11001101100011",
                      17 when "11001101100100",
                      17 when "11001101100101",
                      17 when "11001101100110",
                      17 when "11001101100111",
                      17 when "11001101101000",
                      17 when "11001101101001",
                      17 when "11001101101010",
                      17 when "11001101101011",
                      17 when "11001101101100",
                      17 when "11001101101101",
                      17 when "11001101101110",
                      17 when "11001101101111",
                      17 when "11001101110000",
                      17 when "11001101110001",
                      17 when "11001101110010",
                      17 when "11001101110011",
                      17 when "11001101110100",
                      17 when "11001101110101",
                      17 when "11001101110110",
                      17 when "11001101110111",
                      17 when "11001101111000",
                      17 when "11001101111001",
                      17 when "11001101111010",
                      17 when "11001101111011",
                      17 when "11001101111100",
                      17 when "11001101111101",
                      17 when "11001101111110",
                      17 when "11001101111111",
                      17 when "11001110000000",
                      17 when "11001110000001",
                      17 when "11001110000010",
                      17 when "11001110000011",
                      17 when "11001110000100",
                      17 when "11001110000101",
                      17 when "11001110000110",
                      17 when "11001110000111",
                      17 when "11001110001000",
                      17 when "11001110001001",
                      17 when "11001110001010",
                      17 when "11001110001011",
                      17 when "11001110001100",
                      17 when "11001110001101",
                      17 when "11001110001110",
                      17 when "11001110001111",
                      17 when "11001110010000",
                      17 when "11001110010001",
                      17 when "11001110010010",
                      17 when "11001110010011",
                      17 when "11001110010100",
                      17 when "11001110010101",
                      17 when "11001110010110",
                      17 when "11001110010111",
                      17 when "11001110011000",
                      17 when "11001110011001",
                      17 when "11001110011010",
                      17 when "11001110011011",
                      17 when "11001110011100",
                      17 when "11001110011101",
                      17 when "11001110011110",
                      17 when "11001110011111",
                      17 when "11001110100000",
                      17 when "11001110100001",
                      17 when "11001110100010",
                      17 when "11001110100011",
                      17 when "11001110100100",
                      17 when "11001110100101",
                      17 when "11001110100110",
                      17 when "11001110100111",
                      17 when "11001110101000",
                      17 when "11001110101001",
                      17 when "11001110101010",
                      17 when "11001110101011",
                      17 when "11001110101100",
                      17 when "11001110101101",
                      17 when "11001110101110",
                      17 when "11001110101111",
                      17 when "11001110110000",
                      17 when "11001110110001",
                      17 when "11001110110010",
                      17 when "11001110110011",
                      17 when "11001110110100",
                      17 when "11001110110101",
                      17 when "11001110110110",
                      17 when "11001110110111",
                      17 when "11001110111000",
                      17 when "11001110111001",
                      17 when "11001110111010",
                      17 when "11001110111011",
                      17 when "11001110111100",
                      17 when "11001110111101",
                      17 when "11001110111110",
                      17 when "11001110111111",
                      17 when "11001111000000",
                      17 when "11001111000001",
                      17 when "11001111000010",
                      17 when "11001111000011",
                      17 when "11001111000100",
                      17 when "11001111000101",
                      17 when "11001111000110",
                      17 when "11001111000111",
                      17 when "11001111001000",
                      17 when "11001111001001",
                      17 when "11001111001010",
                      17 when "11001111001011",
                      17 when "11001111001100",
                      17 when "11001111001101",
                      17 when "11001111001110",
                      17 when "11001111001111",
                      17 when "11001111010000",
                      17 when "11001111010001",
                      17 when "11001111010010",
                      17 when "11001111010011",
                      17 when "11001111010100",
                      17 when "11001111010101",
                      17 when "11001111010110",
                      17 when "11001111010111",
                      17 when "11001111011000",
                      17 when "11001111011001",
                      17 when "11001111011010",
                      17 when "11001111011011",
                      17 when "11001111011100",
                      17 when "11001111011101",
                      17 when "11001111011110",
                      17 when "11001111011111",
                      17 when "11001111100000",
                      17 when "11001111100001",
                      17 when "11001111100010",
                      17 when "11001111100011",
                      17 when "11001111100100",
                      17 when "11001111100101",
                      17 when "11001111100110",
                      17 when "11001111100111",
                      17 when "11001111101000",
                      17 when "11001111101001",
                      17 when "11001111101010",
                      17 when "11001111101011",
                      17 when "11001111101100",
                      17 when "11001111101101",
                      17 when "11001111101110",
                      17 when "11001111101111",
                      17 when "11001111110000",
                      17 when "11001111110001",
                      17 when "11001111110010",
                      17 when "11001111110011",
                      17 when "11001111110100",
                      17 when "11001111110101",
                      17 when "11001111110110",
                      17 when "11001111110111",
                      17 when "11001111111000",
                      17 when "11001111111001",
                      17 when "11001111111010",
                      17 when "11001111111011",
                      17 when "11001111111100",
                      17 when "11001111111101",
                      17 when "11001111111110",
                      17 when "11001111111111",
                      17 when "11010000000000",
                      17 when "11010000000001",
                      17 when "11010000000010",
                      17 when "11010000000011",
                      17 when "11010000000100",
                      16 when "11010000000101",
                      16 when "11010000000110",
                      16 when "11010000000111",
                      16 when "11010000001000",
                      16 when "11010000001001",
                      16 when "11010000001010",
                      16 when "11010000001011",
                      16 when "11010000001100",
                      16 when "11010000001101",
                      16 when "11010000001110",
                      16 when "11010000001111",
                      16 when "11010000010000",
                      16 when "11010000010001",
                      16 when "11010000010010",
                      16 when "11010000010011",
                      16 when "11010000010100",
                      16 when "11010000010101",
                      16 when "11010000010110",
                      16 when "11010000010111",
                      16 when "11010000011000",
                      16 when "11010000011001",
                      16 when "11010000011010",
                      16 when "11010000011011",
                      16 when "11010000011100",
                      16 when "11010000011101",
                      16 when "11010000011110",
                      16 when "11010000011111",
                      16 when "11010000100000",
                      16 when "11010000100001",
                      16 when "11010000100010",
                      16 when "11010000100011",
                      16 when "11010000100100",
                      16 when "11010000100101",
                      16 when "11010000100110",
                      16 when "11010000100111",
                      16 when "11010000101000",
                      16 when "11010000101001",
                      16 when "11010000101010",
                      16 when "11010000101011",
                      16 when "11010000101100",
                      16 when "11010000101101",
                      16 when "11010000101110",
                      16 when "11010000101111",
                      16 when "11010000110000",
                      16 when "11010000110001",
                      16 when "11010000110010",
                      16 when "11010000110011",
                      16 when "11010000110100",
                      16 when "11010000110101",
                      16 when "11010000110110",
                      16 when "11010000110111",
                      16 when "11010000111000",
                      16 when "11010000111001",
                      16 when "11010000111010",
                      16 when "11010000111011",
                      16 when "11010000111100",
                      16 when "11010000111101",
                      16 when "11010000111110",
                      16 when "11010000111111",
                      16 when "11010001000000",
                      16 when "11010001000001",
                      16 when "11010001000010",
                      16 when "11010001000011",
                      16 when "11010001000100",
                      16 when "11010001000101",
                      16 when "11010001000110",
                      16 when "11010001000111",
                      16 when "11010001001000",
                      16 when "11010001001001",
                      16 when "11010001001010",
                      16 when "11010001001011",
                      16 when "11010001001100",
                      16 when "11010001001101",
                      16 when "11010001001110",
                      16 when "11010001001111",
                      16 when "11010001010000",
                      16 when "11010001010001",
                      16 when "11010001010010",
                      16 when "11010001010011",
                      16 when "11010001010100",
                      16 when "11010001010101",
                      16 when "11010001010110",
                      16 when "11010001010111",
                      16 when "11010001011000",
                      16 when "11010001011001",
                      16 when "11010001011010",
                      16 when "11010001011011",
                      16 when "11010001011100",
                      16 when "11010001011101",
                      16 when "11010001011110",
                      16 when "11010001011111",
                      16 when "11010001100000",
                      16 when "11010001100001",
                      16 when "11010001100010",
                      16 when "11010001100011",
                      16 when "11010001100100",
                      16 when "11010001100101",
                      16 when "11010001100110",
                      16 when "11010001100111",
                      16 when "11010001101000",
                      16 when "11010001101001",
                      16 when "11010001101010",
                      16 when "11010001101011",
                      16 when "11010001101100",
                      16 when "11010001101101",
                      16 when "11010001101110",
                      16 when "11010001101111",
                      16 when "11010001110000",
                      16 when "11010001110001",
                      16 when "11010001110010",
                      16 when "11010001110011",
                      16 when "11010001110100",
                      16 when "11010001110101",
                      16 when "11010001110110",
                      16 when "11010001110111",
                      16 when "11010001111000",
                      16 when "11010001111001",
                      16 when "11010001111010",
                      16 when "11010001111011",
                      16 when "11010001111100",
                      16 when "11010001111101",
                      16 when "11010001111110",
                      16 when "11010001111111",
                      16 when "11010010000000",
                      16 when "11010010000001",
                      16 when "11010010000010",
                      16 when "11010010000011",
                      16 when "11010010000100",
                      16 when "11010010000101",
                      16 when "11010010000110",
                      16 when "11010010000111",
                      16 when "11010010001000",
                      16 when "11010010001001",
                      16 when "11010010001010",
                      16 when "11010010001011",
                      16 when "11010010001100",
                      16 when "11010010001101",
                      16 when "11010010001110",
                      16 when "11010010001111",
                      16 when "11010010010000",
                      16 when "11010010010001",
                      16 when "11010010010010",
                      16 when "11010010010011",
                      16 when "11010010010100",
                      16 when "11010010010101",
                      16 when "11010010010110",
                      16 when "11010010010111",
                      16 when "11010010011000",
                      16 when "11010010011001",
                      16 when "11010010011010",
                      16 when "11010010011011",
                      16 when "11010010011100",
                      16 when "11010010011101",
                      16 when "11010010011110",
                      16 when "11010010011111",
                      16 when "11010010100000",
                      16 when "11010010100001",
                      16 when "11010010100010",
                      16 when "11010010100011",
                      16 when "11010010100100",
                      16 when "11010010100101",
                      16 when "11010010100110",
                      16 when "11010010100111",
                      16 when "11010010101000",
                      16 when "11010010101001",
                      16 when "11010010101010",
                      16 when "11010010101011",
                      16 when "11010010101100",
                      16 when "11010010101101",
                      16 when "11010010101110",
                      16 when "11010010101111",
                      16 when "11010010110000",
                      16 when "11010010110001",
                      16 when "11010010110010",
                      16 when "11010010110011",
                      16 when "11010010110100",
                      16 when "11010010110101",
                      16 when "11010010110110",
                      16 when "11010010110111",
                      16 when "11010010111000",
                      16 when "11010010111001",
                      16 when "11010010111010",
                      16 when "11010010111011",
                      16 when "11010010111100",
                      16 when "11010010111101",
                      16 when "11010010111110",
                      16 when "11010010111111",
                      16 when "11010011000000",
                      16 when "11010011000001",
                      16 when "11010011000010",
                      16 when "11010011000011",
                      16 when "11010011000100",
                      16 when "11010011000101",
                      16 when "11010011000110",
                      16 when "11010011000111",
                      16 when "11010011001000",
                      16 when "11010011001001",
                      16 when "11010011001010",
                      16 when "11010011001011",
                      16 when "11010011001100",
                      16 when "11010011001101",
                      16 when "11010011001110",
                      16 when "11010011001111",
                      16 when "11010011010000",
                      16 when "11010011010001",
                      16 when "11010011010010",
                      16 when "11010011010011",
                      16 when "11010011010100",
                      16 when "11010011010101",
                      16 when "11010011010110",
                      16 when "11010011010111",
                      16 when "11010011011000",
                      16 when "11010011011001",
                      16 when "11010011011010",
                      16 when "11010011011011",
                      16 when "11010011011100",
                      16 when "11010011011101",
                      16 when "11010011011110",
                      16 when "11010011011111",
                      16 when "11010011100000",
                      16 when "11010011100001",
                      16 when "11010011100010",
                      16 when "11010011100011",
                      16 when "11010011100100",
                      16 when "11010011100101",
                      16 when "11010011100110",
                      16 when "11010011100111",
                      16 when "11010011101000",
                      16 when "11010011101001",
                      16 when "11010011101010",
                      16 when "11010011101011",
                      16 when "11010011101100",
                      16 when "11010011101101",
                      16 when "11010011101110",
                      16 when "11010011101111",
                      16 when "11010011110000",
                      16 when "11010011110001",
                      16 when "11010011110010",
                      16 when "11010011110011",
                      16 when "11010011110100",
                      16 when "11010011110101",
                      16 when "11010011110110",
                      16 when "11010011110111",
                      16 when "11010011111000",
                      16 when "11010011111001",
                      16 when "11010011111010",
                      16 when "11010011111011",
                      16 when "11010011111100",
                      16 when "11010011111101",
                      16 when "11010011111110",
                      16 when "11010011111111",
                      16 when "11010100000000",
                      16 when "11010100000001",
                      16 when "11010100000010",
                      16 when "11010100000011",
                      16 when "11010100000100",
                      16 when "11010100000101",
                      16 when "11010100000110",
                      16 when "11010100000111",
                      16 when "11010100001000",
                      16 when "11010100001001",
                      16 when "11010100001010",
                      16 when "11010100001011",
                      16 when "11010100001100",
                      16 when "11010100001101",
                      16 when "11010100001110",
                      16 when "11010100001111",
                      16 when "11010100010000",
                      16 when "11010100010001",
                      16 when "11010100010010",
                      16 when "11010100010011",
                      16 when "11010100010100",
                      16 when "11010100010101",
                      16 when "11010100010110",
                      16 when "11010100010111",
                      16 when "11010100011000",
                      16 when "11010100011001",
                      16 when "11010100011010",
                      16 when "11010100011011",
                      16 when "11010100011100",
                      16 when "11010100011101",
                      16 when "11010100011110",
                      16 when "11010100011111",
                      16 when "11010100100000",
                      16 when "11010100100001",
                      16 when "11010100100010",
                      16 when "11010100100011",
                      16 when "11010100100100",
                      16 when "11010100100101",
                      16 when "11010100100110",
                      16 when "11010100100111",
                      16 when "11010100101000",
                      16 when "11010100101001",
                      16 when "11010100101010",
                      16 when "11010100101011",
                      16 when "11010100101100",
                      16 when "11010100101101",
                      16 when "11010100101110",
                      16 when "11010100101111",
                      16 when "11010100110000",
                      16 when "11010100110001",
                      16 when "11010100110010",
                      16 when "11010100110011",
                      16 when "11010100110100",
                      16 when "11010100110101",
                      16 when "11010100110110",
                      16 when "11010100110111",
                      16 when "11010100111000",
                      16 when "11010100111001",
                      16 when "11010100111010",
                      16 when "11010100111011",
                      16 when "11010100111100",
                      16 when "11010100111101",
                      16 when "11010100111110",
                      16 when "11010100111111",
                      16 when "11010101000000",
                      16 when "11010101000001",
                      16 when "11010101000010",
                      16 when "11010101000011",
                      16 when "11010101000100",
                      16 when "11010101000101",
                      16 when "11010101000110",
                      16 when "11010101000111",
                      16 when "11010101001000",
                      16 when "11010101001001",
                      16 when "11010101001010",
                      16 when "11010101001011",
                      16 when "11010101001100",
                      16 when "11010101001101",
                      16 when "11010101001110",
                      16 when "11010101001111",
                      16 when "11010101010000",
                      16 when "11010101010001",
                      16 when "11010101010010",
                      16 when "11010101010011",
                      16 when "11010101010100",
                      16 when "11010101010101",
                      16 when "11010101010110",
                      16 when "11010101010111",
                      16 when "11010101011000",
                      16 when "11010101011001",
                      16 when "11010101011010",
                      16 when "11010101011011",
                      16 when "11010101011100",
                      16 when "11010101011101",
                      16 when "11010101011110",
                      16 when "11010101011111",
                      16 when "11010101100000",
                      16 when "11010101100001",
                      16 when "11010101100010",
                      16 when "11010101100011",
                      16 when "11010101100100",
                      16 when "11010101100101",
                      16 when "11010101100110",
                      16 when "11010101100111",
                      16 when "11010101101000",
                      16 when "11010101101001",
                      16 when "11010101101010",
                      16 when "11010101101011",
                      16 when "11010101101100",
                      16 when "11010101101101",
                      16 when "11010101101110",
                      16 when "11010101101111",
                      16 when "11010101110000",
                      16 when "11010101110001",
                      16 when "11010101110010",
                      16 when "11010101110011",
                      16 when "11010101110100",
                      16 when "11010101110101",
                      16 when "11010101110110",
                      16 when "11010101110111",
                      16 when "11010101111000",
                      16 when "11010101111001",
                      16 when "11010101111010",
                      16 when "11010101111011",
                      16 when "11010101111100",
                      16 when "11010101111101",
                      16 when "11010101111110",
                      16 when "11010101111111",
                      16 when "11010110000000",
                      16 when "11010110000001",
                      16 when "11010110000010",
                      16 when "11010110000011",
                      16 when "11010110000100",
                      16 when "11010110000101",
                      16 when "11010110000110",
                      16 when "11010110000111",
                      16 when "11010110001000",
                      16 when "11010110001001",
                      16 when "11010110001010",
                      16 when "11010110001011",
                      16 when "11010110001100",
                      16 when "11010110001101",
                      16 when "11010110001110",
                      16 when "11010110001111",
                      16 when "11010110010000",
                      16 when "11010110010001",
                      16 when "11010110010010",
                      16 when "11010110010011",
                      16 when "11010110010100",
                      16 when "11010110010101",
                      16 when "11010110010110",
                      16 when "11010110010111",
                      16 when "11010110011000",
                      16 when "11010110011001",
                      16 when "11010110011010",
                      16 when "11010110011011",
                      16 when "11010110011100",
                      16 when "11010110011101",
                      16 when "11010110011110",
                      16 when "11010110011111",
                      16 when "11010110100000",
                      16 when "11010110100001",
                      16 when "11010110100010",
                      16 when "11010110100011",
                      16 when "11010110100100",
                      16 when "11010110100101",
                      16 when "11010110100110",
                      16 when "11010110100111",
                      16 when "11010110101000",
                      16 when "11010110101001",
                      16 when "11010110101010",
                      16 when "11010110101011",
                      16 when "11010110101100",
                      16 when "11010110101101",
                      16 when "11010110101110",
                      16 when "11010110101111",
                      16 when "11010110110000",
                      16 when "11010110110001",
                      16 when "11010110110010",
                      16 when "11010110110011",
                      16 when "11010110110100",
                      16 when "11010110110101",
                      16 when "11010110110110",
                      16 when "11010110110111",
                      16 when "11010110111000",
                      16 when "11010110111001",
                      16 when "11010110111010",
                      16 when "11010110111011",
                      16 when "11010110111100",
                      16 when "11010110111101",
                      16 when "11010110111110",
                      16 when "11010110111111",
                      16 when "11010111000000",
                      16 when "11010111000001",
                      16 when "11010111000010",
                      16 when "11010111000011",
                      16 when "11010111000100",
                      16 when "11010111000101",
                      16 when "11010111000110",
                      16 when "11010111000111",
                      16 when "11010111001000",
                      16 when "11010111001001",
                      16 when "11010111001010",
                      16 when "11010111001011",
                      16 when "11010111001100",
                      16 when "11010111001101",
                      16 when "11010111001110",
                      16 when "11010111001111",
                      16 when "11010111010000",
                      16 when "11010111010001",
                      16 when "11010111010010",
                      16 when "11010111010011",
                      16 when "11010111010100",
                      16 when "11010111010101",
                      16 when "11010111010110",
                      16 when "11010111010111",
                      16 when "11010111011000",
                      16 when "11010111011001",
                      16 when "11010111011010",
                      16 when "11010111011011",
                      16 when "11010111011100",
                      16 when "11010111011101",
                      16 when "11010111011110",
                      16 when "11010111011111",
                      16 when "11010111100000",
                      16 when "11010111100001",
                      16 when "11010111100010",
                      16 when "11010111100011",
                      16 when "11010111100100",
                      16 when "11010111100101",
                      16 when "11010111100110",
                      16 when "11010111100111",
                      16 when "11010111101000",
                      16 when "11010111101001",
                      16 when "11010111101010",
                      16 when "11010111101011",
                      16 when "11010111101100",
                      16 when "11010111101101",
                      16 when "11010111101110",
                      16 when "11010111101111",
                      16 when "11010111110000",
                      16 when "11010111110001",
                      16 when "11010111110010",
                      16 when "11010111110011",
                      16 when "11010111110100",
                      16 when "11010111110101",
                      16 when "11010111110110",
                      16 when "11010111110111",
                      16 when "11010111111000",
                      16 when "11010111111001",
                      16 when "11010111111010",
                      16 when "11010111111011",
                      16 when "11010111111100",
                      16 when "11010111111101",
                      16 when "11010111111110",
                      16 when "11010111111111",
                      16 when "11011000000000",
                      16 when "11011000000001",
                      16 when "11011000000010",
                      16 when "11011000000011",
                      16 when "11011000000100",
                      16 when "11011000000101",
                      16 when "11011000000110",
                      16 when "11011000000111",
                      16 when "11011000001000",
                      16 when "11011000001001",
                      16 when "11011000001010",
                      16 when "11011000001011",
                      16 when "11011000001100",
                      16 when "11011000001101",
                      16 when "11011000001110",
                      16 when "11011000001111",
                      16 when "11011000010000",
                      16 when "11011000010001",
                      16 when "11011000010010",
                      16 when "11011000010011",
                      16 when "11011000010100",
                      16 when "11011000010101",
                      16 when "11011000010110",
                      16 when "11011000010111",
                      16 when "11011000011000",
                      16 when "11011000011001",
                      16 when "11011000011010",
                      16 when "11011000011011",
                      16 when "11011000011100",
                      16 when "11011000011101",
                      16 when "11011000011110",
                      16 when "11011000011111",
                      16 when "11011000100000",
                      16 when "11011000100001",
                      16 when "11011000100010",
                      16 when "11011000100011",
                      16 when "11011000100100",
                      16 when "11011000100101",
                      16 when "11011000100110",
                      16 when "11011000100111",
                      16 when "11011000101000",
                      16 when "11011000101001",
                      16 when "11011000101010",
                      16 when "11011000101011",
                      16 when "11011000101100",
                      16 when "11011000101101",
                      16 when "11011000101110",
                      16 when "11011000101111",
                      16 when "11011000110000",
                      16 when "11011000110001",
                      16 when "11011000110010",
                      16 when "11011000110011",
                      16 when "11011000110100",
                      16 when "11011000110101",
                      16 when "11011000110110",
                      16 when "11011000110111",
                      16 when "11011000111000",
                      16 when "11011000111001",
                      16 when "11011000111010",
                      16 when "11011000111011",
                      16 when "11011000111100",
                      16 when "11011000111101",
                      16 when "11011000111110",
                      16 when "11011000111111",
                      16 when "11011001000000",
                      16 when "11011001000001",
                      16 when "11011001000010",
                      16 when "11011001000011",
                      16 when "11011001000100",
                      16 when "11011001000101",
                      16 when "11011001000110",
                      16 when "11011001000111",
                      16 when "11011001001000",
                      16 when "11011001001001",
                      16 when "11011001001010",
                      16 when "11011001001011",
                      16 when "11011001001100",
                      16 when "11011001001101",
                      16 when "11011001001110",
                      16 when "11011001001111",
                      16 when "11011001010000",
                      16 when "11011001010001",
                      16 when "11011001010010",
                      16 when "11011001010011",
                      16 when "11011001010100",
                      16 when "11011001010101",
                      16 when "11011001010110",
                      16 when "11011001010111",
                      16 when "11011001011000",
                      16 when "11011001011001",
                      16 when "11011001011010",
                      16 when "11011001011011",
                      16 when "11011001011100",
                      16 when "11011001011101",
                      16 when "11011001011110",
                      16 when "11011001011111",
                      16 when "11011001100000",
                      16 when "11011001100001",
                      16 when "11011001100010",
                      16 when "11011001100011",
                      16 when "11011001100100",
                      16 when "11011001100101",
                      16 when "11011001100110",
                      16 when "11011001100111",
                      16 when "11011001101000",
                      16 when "11011001101001",
                      16 when "11011001101010",
                      16 when "11011001101011",
                      16 when "11011001101100",
                      16 when "11011001101101",
                      16 when "11011001101110",
                      16 when "11011001101111",
                      16 when "11011001110000",
                      16 when "11011001110001",
                      16 when "11011001110010",
                      16 when "11011001110011",
                      16 when "11011001110100",
                      16 when "11011001110101",
                      16 when "11011001110110",
                      16 when "11011001110111",
                      16 when "11011001111000",
                      16 when "11011001111001",
                      16 when "11011001111010",
                      16 when "11011001111011",
                      16 when "11011001111100",
                      16 when "11011001111101",
                      16 when "11011001111110",
                      16 when "11011001111111",
                      16 when "11011010000000",
                      16 when "11011010000001",
                      16 when "11011010000010",
                      16 when "11011010000011",
                      16 when "11011010000100",
                      16 when "11011010000101",
                      16 when "11011010000110",
                      16 when "11011010000111",
                      16 when "11011010001000",
                      16 when "11011010001001",
                      16 when "11011010001010",
                      16 when "11011010001011",
                      16 when "11011010001100",
                      16 when "11011010001101",
                      16 when "11011010001110",
                      16 when "11011010001111",
                      16 when "11011010010000",
                      16 when "11011010010001",
                      16 when "11011010010010",
                      16 when "11011010010011",
                      16 when "11011010010100",
                      16 when "11011010010101",
                      16 when "11011010010110",
                      16 when "11011010010111",
                      16 when "11011010011000",
                      16 when "11011010011001",
                      16 when "11011010011010",
                      16 when "11011010011011",
                      16 when "11011010011100",
                      16 when "11011010011101",
                      16 when "11011010011110",
                      16 when "11011010011111",
                      16 when "11011010100000",
                      16 when "11011010100001",
                      16 when "11011010100010",
                      16 when "11011010100011",
                      16 when "11011010100100",
                      16 when "11011010100101",
                      16 when "11011010100110",
                      16 when "11011010100111",
                      16 when "11011010101000",
                      16 when "11011010101001",
                      16 when "11011010101010",
                      16 when "11011010101011",
                      16 when "11011010101100",
                      16 when "11011010101101",
                      16 when "11011010101110",
                      16 when "11011010101111",
                      16 when "11011010110000",
                      16 when "11011010110001",
                      16 when "11011010110010",
                      16 when "11011010110011",
                      16 when "11011010110100",
                      16 when "11011010110101",
                      16 when "11011010110110",
                      16 when "11011010110111",
                      16 when "11011010111000",
                      16 when "11011010111001",
                      16 when "11011010111010",
                      16 when "11011010111011",
                      16 when "11011010111100",
                      16 when "11011010111101",
                      16 when "11011010111110",
                      16 when "11011010111111",
                      16 when "11011011000000",
                      16 when "11011011000001",
                      16 when "11011011000010",
                      16 when "11011011000011",
                      16 when "11011011000100",
                      16 when "11011011000101",
                      16 when "11011011000110",
                      16 when "11011011000111",
                      16 when "11011011001000",
                      16 when "11011011001001",
                      16 when "11011011001010",
                      16 when "11011011001011",
                      16 when "11011011001100",
                      16 when "11011011001101",
                      16 when "11011011001110",
                      16 when "11011011001111",
                      16 when "11011011010000",
                      16 when "11011011010001",
                      16 when "11011011010010",
                      16 when "11011011010011",
                      16 when "11011011010100",
                      16 when "11011011010101",
                      16 when "11011011010110",
                      16 when "11011011010111",
                      16 when "11011011011000",
                      16 when "11011011011001",
                      16 when "11011011011010",
                      16 when "11011011011011",
                      16 when "11011011011100",
                      16 when "11011011011101",
                      16 when "11011011011110",
                      16 when "11011011011111",
                      16 when "11011011100000",
                      16 when "11011011100001",
                      16 when "11011011100010",
                      16 when "11011011100011",
                      16 when "11011011100100",
                      16 when "11011011100101",
                      16 when "11011011100110",
                      16 when "11011011100111",
                      16 when "11011011101000",
                      16 when "11011011101001",
                      16 when "11011011101010",
                      16 when "11011011101011",
                      16 when "11011011101100",
                      16 when "11011011101101",
                      16 when "11011011101110",
                      16 when "11011011101111",
                      16 when "11011011110000",
                      16 when "11011011110001",
                      16 when "11011011110010",
                      16 when "11011011110011",
                      16 when "11011011110100",
                      16 when "11011011110101",
                      16 when "11011011110110",
                      16 when "11011011110111",
                      16 when "11011011111000",
                      16 when "11011011111001",
                      16 when "11011011111010",
                      16 when "11011011111011",
                      16 when "11011011111100",
                      16 when "11011011111101",
                      16 when "11011011111110",
                      16 when "11011011111111",
                      16 when "11011100000000",
                      16 when "11011100000001",
                      16 when "11011100000010",
                      16 when "11011100000011",
                      16 when "11011100000100",
                      16 when "11011100000101",
                      16 when "11011100000110",
                      16 when "11011100000111",
                      16 when "11011100001000",
                      16 when "11011100001001",
                      16 when "11011100001010",
                      16 when "11011100001011",
                      16 when "11011100001100",
                      16 when "11011100001101",
                      16 when "11011100001110",
                      16 when "11011100001111",
                      16 when "11011100010000",
                      16 when "11011100010001",
                      16 when "11011100010010",
                      16 when "11011100010011",
                      16 when "11011100010100",
                      16 when "11011100010101",
                      16 when "11011100010110",
                      16 when "11011100010111",
                      16 when "11011100011000",
                      16 when "11011100011001",
                      16 when "11011100011010",
                      16 when "11011100011011",
                      16 when "11011100011100",
                      16 when "11011100011101",
                      16 when "11011100011110",
                      16 when "11011100011111",
                      16 when "11011100100000",
                      16 when "11011100100001",
                      16 when "11011100100010",
                      16 when "11011100100011",
                      16 when "11011100100100",
                      16 when "11011100100101",
                      16 when "11011100100110",
                      16 when "11011100100111",
                      16 when "11011100101000",
                      16 when "11011100101001",
                      16 when "11011100101010",
                      16 when "11011100101011",
                      16 when "11011100101100",
                      16 when "11011100101101",
                      16 when "11011100101110",
                      16 when "11011100101111",
                      16 when "11011100110000",
                      16 when "11011100110001",
                      16 when "11011100110010",
                      16 when "11011100110011",
                      16 when "11011100110100",
                      16 when "11011100110101",
                      16 when "11011100110110",
                      16 when "11011100110111",
                      16 when "11011100111000",
                      16 when "11011100111001",
                      16 when "11011100111010",
                      16 when "11011100111011",
                      16 when "11011100111100",
                      16 when "11011100111101",
                      16 when "11011100111110",
                      16 when "11011100111111",
                      16 when "11011101000000",
                      16 when "11011101000001",
                      16 when "11011101000010",
                      16 when "11011101000011",
                      16 when "11011101000100",
                      16 when "11011101000101",
                      16 when "11011101000110",
                      16 when "11011101000111",
                      16 when "11011101001000",
                      16 when "11011101001001",
                      16 when "11011101001010",
                      16 when "11011101001011",
                      16 when "11011101001100",
                      16 when "11011101001101",
                      16 when "11011101001110",
                      16 when "11011101001111",
                      16 when "11011101010000",
                      16 when "11011101010001",
                      16 when "11011101010010",
                      16 when "11011101010011",
                      16 when "11011101010100",
                      16 when "11011101010101",
                      16 when "11011101010110",
                      16 when "11011101010111",
                      16 when "11011101011000",
                      16 when "11011101011001",
                      16 when "11011101011010",
                      16 when "11011101011011",
                      16 when "11011101011100",
                      16 when "11011101011101",
                      16 when "11011101011110",
                      16 when "11011101011111",
                      15 when "11011101100000",
                      15 when "11011101100001",
                      15 when "11011101100010",
                      15 when "11011101100011",
                      15 when "11011101100100",
                      15 when "11011101100101",
                      15 when "11011101100110",
                      15 when "11011101100111",
                      15 when "11011101101000",
                      15 when "11011101101001",
                      15 when "11011101101010",
                      15 when "11011101101011",
                      15 when "11011101101100",
                      15 when "11011101101101",
                      15 when "11011101101110",
                      15 when "11011101101111",
                      15 when "11011101110000",
                      15 when "11011101110001",
                      15 when "11011101110010",
                      15 when "11011101110011",
                      15 when "11011101110100",
                      15 when "11011101110101",
                      15 when "11011101110110",
                      15 when "11011101110111",
                      15 when "11011101111000",
                      15 when "11011101111001",
                      15 when "11011101111010",
                      15 when "11011101111011",
                      15 when "11011101111100",
                      15 when "11011101111101",
                      15 when "11011101111110",
                      15 when "11011101111111",
                      15 when "11011110000000",
                      15 when "11011110000001",
                      15 when "11011110000010",
                      15 when "11011110000011",
                      15 when "11011110000100",
                      15 when "11011110000101",
                      15 when "11011110000110",
                      15 when "11011110000111",
                      15 when "11011110001000",
                      15 when "11011110001001",
                      15 when "11011110001010",
                      15 when "11011110001011",
                      15 when "11011110001100",
                      15 when "11011110001101",
                      15 when "11011110001110",
                      15 when "11011110001111",
                      15 when "11011110010000",
                      15 when "11011110010001",
                      15 when "11011110010010",
                      15 when "11011110010011",
                      15 when "11011110010100",
                      15 when "11011110010101",
                      15 when "11011110010110",
                      15 when "11011110010111",
                      15 when "11011110011000",
                      15 when "11011110011001",
                      15 when "11011110011010",
                      15 when "11011110011011",
                      15 when "11011110011100",
                      15 when "11011110011101",
                      15 when "11011110011110",
                      15 when "11011110011111",
                      15 when "11011110100000",
                      15 when "11011110100001",
                      15 when "11011110100010",
                      15 when "11011110100011",
                      15 when "11011110100100",
                      15 when "11011110100101",
                      15 when "11011110100110",
                      15 when "11011110100111",
                      15 when "11011110101000",
                      15 when "11011110101001",
                      15 when "11011110101010",
                      15 when "11011110101011",
                      15 when "11011110101100",
                      15 when "11011110101101",
                      15 when "11011110101110",
                      15 when "11011110101111",
                      15 when "11011110110000",
                      15 when "11011110110001",
                      15 when "11011110110010",
                      15 when "11011110110011",
                      15 when "11011110110100",
                      15 when "11011110110101",
                      15 when "11011110110110",
                      15 when "11011110110111",
                      15 when "11011110111000",
                      15 when "11011110111001",
                      15 when "11011110111010",
                      15 when "11011110111011",
                      15 when "11011110111100",
                      15 when "11011110111101",
                      15 when "11011110111110",
                      15 when "11011110111111",
                      15 when "11011111000000",
                      15 when "11011111000001",
                      15 when "11011111000010",
                      15 when "11011111000011",
                      15 when "11011111000100",
                      15 when "11011111000101",
                      15 when "11011111000110",
                      15 when "11011111000111",
                      15 when "11011111001000",
                      15 when "11011111001001",
                      15 when "11011111001010",
                      15 when "11011111001011",
                      15 when "11011111001100",
                      15 when "11011111001101",
                      15 when "11011111001110",
                      15 when "11011111001111",
                      15 when "11011111010000",
                      15 when "11011111010001",
                      15 when "11011111010010",
                      15 when "11011111010011",
                      15 when "11011111010100",
                      15 when "11011111010101",
                      15 when "11011111010110",
                      15 when "11011111010111",
                      15 when "11011111011000",
                      15 when "11011111011001",
                      15 when "11011111011010",
                      15 when "11011111011011",
                      15 when "11011111011100",
                      15 when "11011111011101",
                      15 when "11011111011110",
                      15 when "11011111011111",
                      15 when "11011111100000",
                      15 when "11011111100001",
                      15 when "11011111100010",
                      15 when "11011111100011",
                      15 when "11011111100100",
                      15 when "11011111100101",
                      15 when "11011111100110",
                      15 when "11011111100111",
                      15 when "11011111101000",
                      15 when "11011111101001",
                      15 when "11011111101010",
                      15 when "11011111101011",
                      15 when "11011111101100",
                      15 when "11011111101101",
                      15 when "11011111101110",
                      15 when "11011111101111",
                      15 when "11011111110000",
                      15 when "11011111110001",
                      15 when "11011111110010",
                      15 when "11011111110011",
                      15 when "11011111110100",
                      15 when "11011111110101",
                      15 when "11011111110110",
                      15 when "11011111110111",
                      15 when "11011111111000",
                      15 when "11011111111001",
                      15 when "11011111111010",
                      15 when "11011111111011",
                      15 when "11011111111100",
                      15 when "11011111111101",
                      15 when "11011111111110",
                      15 when "11011111111111",
                      15 when "11100000000000",
                      15 when "11100000000001",
                      15 when "11100000000010",
                      15 when "11100000000011",
                      15 when "11100000000100",
                      15 when "11100000000101",
                      15 when "11100000000110",
                      15 when "11100000000111",
                      15 when "11100000001000",
                      15 when "11100000001001",
                      15 when "11100000001010",
                      15 when "11100000001011",
                      15 when "11100000001100",
                      15 when "11100000001101",
                      15 when "11100000001110",
                      15 when "11100000001111",
                      15 when "11100000010000",
                      15 when "11100000010001",
                      15 when "11100000010010",
                      15 when "11100000010011",
                      15 when "11100000010100",
                      15 when "11100000010101",
                      15 when "11100000010110",
                      15 when "11100000010111",
                      15 when "11100000011000",
                      15 when "11100000011001",
                      15 when "11100000011010",
                      15 when "11100000011011",
                      15 when "11100000011100",
                      15 when "11100000011101",
                      15 when "11100000011110",
                      15 when "11100000011111",
                      15 when "11100000100000",
                      15 when "11100000100001",
                      15 when "11100000100010",
                      15 when "11100000100011",
                      15 when "11100000100100",
                      15 when "11100000100101",
                      15 when "11100000100110",
                      15 when "11100000100111",
                      15 when "11100000101000",
                      15 when "11100000101001",
                      15 when "11100000101010",
                      15 when "11100000101011",
                      15 when "11100000101100",
                      15 when "11100000101101",
                      15 when "11100000101110",
                      15 when "11100000101111",
                      15 when "11100000110000",
                      15 when "11100000110001",
                      15 when "11100000110010",
                      15 when "11100000110011",
                      15 when "11100000110100",
                      15 when "11100000110101",
                      15 when "11100000110110",
                      15 when "11100000110111",
                      15 when "11100000111000",
                      15 when "11100000111001",
                      15 when "11100000111010",
                      15 when "11100000111011",
                      15 when "11100000111100",
                      15 when "11100000111101",
                      15 when "11100000111110",
                      15 when "11100000111111",
                      15 when "11100001000000",
                      15 when "11100001000001",
                      15 when "11100001000010",
                      15 when "11100001000011",
                      15 when "11100001000100",
                      15 when "11100001000101",
                      15 when "11100001000110",
                      15 when "11100001000111",
                      15 when "11100001001000",
                      15 when "11100001001001",
                      15 when "11100001001010",
                      15 when "11100001001011",
                      15 when "11100001001100",
                      15 when "11100001001101",
                      15 when "11100001001110",
                      15 when "11100001001111",
                      15 when "11100001010000",
                      15 when "11100001010001",
                      15 when "11100001010010",
                      15 when "11100001010011",
                      15 when "11100001010100",
                      15 when "11100001010101",
                      15 when "11100001010110",
                      15 when "11100001010111",
                      15 when "11100001011000",
                      15 when "11100001011001",
                      15 when "11100001011010",
                      15 when "11100001011011",
                      15 when "11100001011100",
                      15 when "11100001011101",
                      15 when "11100001011110",
                      15 when "11100001011111",
                      15 when "11100001100000",
                      15 when "11100001100001",
                      15 when "11100001100010",
                      15 when "11100001100011",
                      15 when "11100001100100",
                      15 when "11100001100101",
                      15 when "11100001100110",
                      15 when "11100001100111",
                      15 when "11100001101000",
                      15 when "11100001101001",
                      15 when "11100001101010",
                      15 when "11100001101011",
                      15 when "11100001101100",
                      15 when "11100001101101",
                      15 when "11100001101110",
                      15 when "11100001101111",
                      15 when "11100001110000",
                      15 when "11100001110001",
                      15 when "11100001110010",
                      15 when "11100001110011",
                      15 when "11100001110100",
                      15 when "11100001110101",
                      15 when "11100001110110",
                      15 when "11100001110111",
                      15 when "11100001111000",
                      15 when "11100001111001",
                      15 when "11100001111010",
                      15 when "11100001111011",
                      15 when "11100001111100",
                      15 when "11100001111101",
                      15 when "11100001111110",
                      15 when "11100001111111",
                      15 when "11100010000000",
                      15 when "11100010000001",
                      15 when "11100010000010",
                      15 when "11100010000011",
                      15 when "11100010000100",
                      15 when "11100010000101",
                      15 when "11100010000110",
                      15 when "11100010000111",
                      15 when "11100010001000",
                      15 when "11100010001001",
                      15 when "11100010001010",
                      15 when "11100010001011",
                      15 when "11100010001100",
                      15 when "11100010001101",
                      15 when "11100010001110",
                      15 when "11100010001111",
                      15 when "11100010010000",
                      15 when "11100010010001",
                      15 when "11100010010010",
                      15 when "11100010010011",
                      15 when "11100010010100",
                      15 when "11100010010101",
                      15 when "11100010010110",
                      15 when "11100010010111",
                      15 when "11100010011000",
                      15 when "11100010011001",
                      15 when "11100010011010",
                      15 when "11100010011011",
                      15 when "11100010011100",
                      15 when "11100010011101",
                      15 when "11100010011110",
                      15 when "11100010011111",
                      15 when "11100010100000",
                      15 when "11100010100001",
                      15 when "11100010100010",
                      15 when "11100010100011",
                      15 when "11100010100100",
                      15 when "11100010100101",
                      15 when "11100010100110",
                      15 when "11100010100111",
                      15 when "11100010101000",
                      15 when "11100010101001",
                      15 when "11100010101010",
                      15 when "11100010101011",
                      15 when "11100010101100",
                      15 when "11100010101101",
                      15 when "11100010101110",
                      15 when "11100010101111",
                      15 when "11100010110000",
                      15 when "11100010110001",
                      15 when "11100010110010",
                      15 when "11100010110011",
                      15 when "11100010110100",
                      15 when "11100010110101",
                      15 when "11100010110110",
                      15 when "11100010110111",
                      15 when "11100010111000",
                      15 when "11100010111001",
                      15 when "11100010111010",
                      15 when "11100010111011",
                      15 when "11100010111100",
                      15 when "11100010111101",
                      15 when "11100010111110",
                      15 when "11100010111111",
                      15 when "11100011000000",
                      15 when "11100011000001",
                      15 when "11100011000010",
                      15 when "11100011000011",
                      15 when "11100011000100",
                      15 when "11100011000101",
                      15 when "11100011000110",
                      15 when "11100011000111",
                      15 when "11100011001000",
                      15 when "11100011001001",
                      15 when "11100011001010",
                      15 when "11100011001011",
                      15 when "11100011001100",
                      15 when "11100011001101",
                      15 when "11100011001110",
                      15 when "11100011001111",
                      15 when "11100011010000",
                      15 when "11100011010001",
                      15 when "11100011010010",
                      15 when "11100011010011",
                      15 when "11100011010100",
                      15 when "11100011010101",
                      15 when "11100011010110",
                      15 when "11100011010111",
                      15 when "11100011011000",
                      15 when "11100011011001",
                      15 when "11100011011010",
                      15 when "11100011011011",
                      15 when "11100011011100",
                      15 when "11100011011101",
                      15 when "11100011011110",
                      15 when "11100011011111",
                      15 when "11100011100000",
                      15 when "11100011100001",
                      15 when "11100011100010",
                      15 when "11100011100011",
                      15 when "11100011100100",
                      15 when "11100011100101",
                      15 when "11100011100110",
                      15 when "11100011100111",
                      15 when "11100011101000",
                      15 when "11100011101001",
                      15 when "11100011101010",
                      15 when "11100011101011",
                      15 when "11100011101100",
                      15 when "11100011101101",
                      15 when "11100011101110",
                      15 when "11100011101111",
                      15 when "11100011110000",
                      15 when "11100011110001",
                      15 when "11100011110010",
                      15 when "11100011110011",
                      15 when "11100011110100",
                      15 when "11100011110101",
                      15 when "11100011110110",
                      15 when "11100011110111",
                      15 when "11100011111000",
                      15 when "11100011111001",
                      15 when "11100011111010",
                      15 when "11100011111011",
                      15 when "11100011111100",
                      15 when "11100011111101",
                      15 when "11100011111110",
                      15 when "11100011111111",
                      15 when "11100100000000",
                      15 when "11100100000001",
                      15 when "11100100000010",
                      15 when "11100100000011",
                      15 when "11100100000100",
                      15 when "11100100000101",
                      15 when "11100100000110",
                      15 when "11100100000111",
                      15 when "11100100001000",
                      15 when "11100100001001",
                      15 when "11100100001010",
                      15 when "11100100001011",
                      15 when "11100100001100",
                      15 when "11100100001101",
                      15 when "11100100001110",
                      15 when "11100100001111",
                      15 when "11100100010000",
                      15 when "11100100010001",
                      15 when "11100100010010",
                      15 when "11100100010011",
                      15 when "11100100010100",
                      15 when "11100100010101",
                      15 when "11100100010110",
                      15 when "11100100010111",
                      15 when "11100100011000",
                      15 when "11100100011001",
                      15 when "11100100011010",
                      15 when "11100100011011",
                      15 when "11100100011100",
                      15 when "11100100011101",
                      15 when "11100100011110",
                      15 when "11100100011111",
                      15 when "11100100100000",
                      15 when "11100100100001",
                      15 when "11100100100010",
                      15 when "11100100100011",
                      15 when "11100100100100",
                      15 when "11100100100101",
                      15 when "11100100100110",
                      15 when "11100100100111",
                      15 when "11100100101000",
                      15 when "11100100101001",
                      15 when "11100100101010",
                      15 when "11100100101011",
                      15 when "11100100101100",
                      15 when "11100100101101",
                      15 when "11100100101110",
                      15 when "11100100101111",
                      15 when "11100100110000",
                      15 when "11100100110001",
                      15 when "11100100110010",
                      15 when "11100100110011",
                      15 when "11100100110100",
                      15 when "11100100110101",
                      15 when "11100100110110",
                      15 when "11100100110111",
                      15 when "11100100111000",
                      15 when "11100100111001",
                      15 when "11100100111010",
                      15 when "11100100111011",
                      15 when "11100100111100",
                      15 when "11100100111101",
                      15 when "11100100111110",
                      15 when "11100100111111",
                      15 when "11100101000000",
                      15 when "11100101000001",
                      15 when "11100101000010",
                      15 when "11100101000011",
                      15 when "11100101000100",
                      15 when "11100101000101",
                      15 when "11100101000110",
                      15 when "11100101000111",
                      15 when "11100101001000",
                      15 when "11100101001001",
                      15 when "11100101001010",
                      15 when "11100101001011",
                      15 when "11100101001100",
                      15 when "11100101001101",
                      15 when "11100101001110",
                      15 when "11100101001111",
                      15 when "11100101010000",
                      15 when "11100101010001",
                      15 when "11100101010010",
                      15 when "11100101010011",
                      15 when "11100101010100",
                      15 when "11100101010101",
                      15 when "11100101010110",
                      15 when "11100101010111",
                      15 when "11100101011000",
                      15 when "11100101011001",
                      15 when "11100101011010",
                      15 when "11100101011011",
                      15 when "11100101011100",
                      15 when "11100101011101",
                      15 when "11100101011110",
                      15 when "11100101011111",
                      15 when "11100101100000",
                      15 when "11100101100001",
                      15 when "11100101100010",
                      15 when "11100101100011",
                      15 when "11100101100100",
                      15 when "11100101100101",
                      15 when "11100101100110",
                      15 when "11100101100111",
                      15 when "11100101101000",
                      15 when "11100101101001",
                      15 when "11100101101010",
                      15 when "11100101101011",
                      15 when "11100101101100",
                      15 when "11100101101101",
                      15 when "11100101101110",
                      15 when "11100101101111",
                      15 when "11100101110000",
                      15 when "11100101110001",
                      15 when "11100101110010",
                      15 when "11100101110011",
                      15 when "11100101110100",
                      15 when "11100101110101",
                      15 when "11100101110110",
                      15 when "11100101110111",
                      15 when "11100101111000",
                      15 when "11100101111001",
                      15 when "11100101111010",
                      15 when "11100101111011",
                      15 when "11100101111100",
                      15 when "11100101111101",
                      15 when "11100101111110",
                      15 when "11100101111111",
                      15 when "11100110000000",
                      15 when "11100110000001",
                      15 when "11100110000010",
                      15 when "11100110000011",
                      15 when "11100110000100",
                      15 when "11100110000101",
                      15 when "11100110000110",
                      15 when "11100110000111",
                      15 when "11100110001000",
                      15 when "11100110001001",
                      15 when "11100110001010",
                      15 when "11100110001011",
                      15 when "11100110001100",
                      15 when "11100110001101",
                      15 when "11100110001110",
                      15 when "11100110001111",
                      15 when "11100110010000",
                      15 when "11100110010001",
                      15 when "11100110010010",
                      15 when "11100110010011",
                      15 when "11100110010100",
                      15 when "11100110010101",
                      15 when "11100110010110",
                      15 when "11100110010111",
                      15 when "11100110011000",
                      15 when "11100110011001",
                      15 when "11100110011010",
                      15 when "11100110011011",
                      15 when "11100110011100",
                      15 when "11100110011101",
                      15 when "11100110011110",
                      15 when "11100110011111",
                      15 when "11100110100000",
                      15 when "11100110100001",
                      15 when "11100110100010",
                      15 when "11100110100011",
                      15 when "11100110100100",
                      15 when "11100110100101",
                      15 when "11100110100110",
                      15 when "11100110100111",
                      15 when "11100110101000",
                      15 when "11100110101001",
                      15 when "11100110101010",
                      15 when "11100110101011",
                      15 when "11100110101100",
                      15 when "11100110101101",
                      15 when "11100110101110",
                      15 when "11100110101111",
                      15 when "11100110110000",
                      15 when "11100110110001",
                      15 when "11100110110010",
                      15 when "11100110110011",
                      15 when "11100110110100",
                      15 when "11100110110101",
                      15 when "11100110110110",
                      15 when "11100110110111",
                      15 when "11100110111000",
                      15 when "11100110111001",
                      15 when "11100110111010",
                      15 when "11100110111011",
                      15 when "11100110111100",
                      15 when "11100110111101",
                      15 when "11100110111110",
                      15 when "11100110111111",
                      15 when "11100111000000",
                      15 when "11100111000001",
                      15 when "11100111000010",
                      15 when "11100111000011",
                      15 when "11100111000100",
                      15 when "11100111000101",
                      15 when "11100111000110",
                      15 when "11100111000111",
                      15 when "11100111001000",
                      15 when "11100111001001",
                      15 when "11100111001010",
                      15 when "11100111001011",
                      15 when "11100111001100",
                      15 when "11100111001101",
                      15 when "11100111001110",
                      15 when "11100111001111",
                      15 when "11100111010000",
                      15 when "11100111010001",
                      15 when "11100111010010",
                      15 when "11100111010011",
                      15 when "11100111010100",
                      15 when "11100111010101",
                      15 when "11100111010110",
                      15 when "11100111010111",
                      15 when "11100111011000",
                      15 when "11100111011001",
                      15 when "11100111011010",
                      15 when "11100111011011",
                      15 when "11100111011100",
                      15 when "11100111011101",
                      15 when "11100111011110",
                      15 when "11100111011111",
                      15 when "11100111100000",
                      15 when "11100111100001",
                      15 when "11100111100010",
                      15 when "11100111100011",
                      15 when "11100111100100",
                      15 when "11100111100101",
                      15 when "11100111100110",
                      15 when "11100111100111",
                      15 when "11100111101000",
                      15 when "11100111101001",
                      15 when "11100111101010",
                      15 when "11100111101011",
                      15 when "11100111101100",
                      15 when "11100111101101",
                      15 when "11100111101110",
                      15 when "11100111101111",
                      15 when "11100111110000",
                      15 when "11100111110001",
                      15 when "11100111110010",
                      15 when "11100111110011",
                      15 when "11100111110100",
                      15 when "11100111110101",
                      15 when "11100111110110",
                      15 when "11100111110111",
                      15 when "11100111111000",
                      15 when "11100111111001",
                      15 when "11100111111010",
                      15 when "11100111111011",
                      15 when "11100111111100",
                      15 when "11100111111101",
                      15 when "11100111111110",
                      15 when "11100111111111",
                      15 when "11101000000000",
                      15 when "11101000000001",
                      15 when "11101000000010",
                      15 when "11101000000011",
                      15 when "11101000000100",
                      15 when "11101000000101",
                      15 when "11101000000110",
                      15 when "11101000000111",
                      15 when "11101000001000",
                      15 when "11101000001001",
                      15 when "11101000001010",
                      15 when "11101000001011",
                      15 when "11101000001100",
                      15 when "11101000001101",
                      15 when "11101000001110",
                      15 when "11101000001111",
                      15 when "11101000010000",
                      15 when "11101000010001",
                      15 when "11101000010010",
                      15 when "11101000010011",
                      15 when "11101000010100",
                      15 when "11101000010101",
                      15 when "11101000010110",
                      15 when "11101000010111",
                      15 when "11101000011000",
                      15 when "11101000011001",
                      15 when "11101000011010",
                      15 when "11101000011011",
                      15 when "11101000011100",
                      15 when "11101000011101",
                      15 when "11101000011110",
                      15 when "11101000011111",
                      15 when "11101000100000",
                      15 when "11101000100001",
                      15 when "11101000100010",
                      15 when "11101000100011",
                      15 when "11101000100100",
                      15 when "11101000100101",
                      15 when "11101000100110",
                      15 when "11101000100111",
                      15 when "11101000101000",
                      15 when "11101000101001",
                      15 when "11101000101010",
                      15 when "11101000101011",
                      15 when "11101000101100",
                      15 when "11101000101101",
                      15 when "11101000101110",
                      15 when "11101000101111",
                      15 when "11101000110000",
                      15 when "11101000110001",
                      15 when "11101000110010",
                      15 when "11101000110011",
                      15 when "11101000110100",
                      15 when "11101000110101",
                      15 when "11101000110110",
                      15 when "11101000110111",
                      15 when "11101000111000",
                      15 when "11101000111001",
                      15 when "11101000111010",
                      15 when "11101000111011",
                      15 when "11101000111100",
                      15 when "11101000111101",
                      15 when "11101000111110",
                      15 when "11101000111111",
                      15 when "11101001000000",
                      15 when "11101001000001",
                      15 when "11101001000010",
                      15 when "11101001000011",
                      15 when "11101001000100",
                      15 when "11101001000101",
                      15 when "11101001000110",
                      15 when "11101001000111",
                      15 when "11101001001000",
                      15 when "11101001001001",
                      15 when "11101001001010",
                      15 when "11101001001011",
                      15 when "11101001001100",
                      15 when "11101001001101",
                      15 when "11101001001110",
                      15 when "11101001001111",
                      15 when "11101001010000",
                      15 when "11101001010001",
                      15 when "11101001010010",
                      15 when "11101001010011",
                      15 when "11101001010100",
                      15 when "11101001010101",
                      15 when "11101001010110",
                      15 when "11101001010111",
                      15 when "11101001011000",
                      15 when "11101001011001",
                      15 when "11101001011010",
                      15 when "11101001011011",
                      15 when "11101001011100",
                      15 when "11101001011101",
                      15 when "11101001011110",
                      15 when "11101001011111",
                      15 when "11101001100000",
                      15 when "11101001100001",
                      15 when "11101001100010",
                      15 when "11101001100011",
                      15 when "11101001100100",
                      15 when "11101001100101",
                      15 when "11101001100110",
                      15 when "11101001100111",
                      15 when "11101001101000",
                      15 when "11101001101001",
                      15 when "11101001101010",
                      15 when "11101001101011",
                      15 when "11101001101100",
                      15 when "11101001101101",
                      15 when "11101001101110",
                      15 when "11101001101111",
                      15 when "11101001110000",
                      15 when "11101001110001",
                      15 when "11101001110010",
                      15 when "11101001110011",
                      15 when "11101001110100",
                      15 when "11101001110101",
                      15 when "11101001110110",
                      15 when "11101001110111",
                      15 when "11101001111000",
                      15 when "11101001111001",
                      15 when "11101001111010",
                      15 when "11101001111011",
                      15 when "11101001111100",
                      15 when "11101001111101",
                      15 when "11101001111110",
                      15 when "11101001111111",
                      15 when "11101010000000",
                      15 when "11101010000001",
                      15 when "11101010000010",
                      15 when "11101010000011",
                      15 when "11101010000100",
                      15 when "11101010000101",
                      15 when "11101010000110",
                      15 when "11101010000111",
                      15 when "11101010001000",
                      15 when "11101010001001",
                      15 when "11101010001010",
                      15 when "11101010001011",
                      15 when "11101010001100",
                      15 when "11101010001101",
                      15 when "11101010001110",
                      15 when "11101010001111",
                      15 when "11101010010000",
                      15 when "11101010010001",
                      15 when "11101010010010",
                      15 when "11101010010011",
                      15 when "11101010010100",
                      15 when "11101010010101",
                      15 when "11101010010110",
                      15 when "11101010010111",
                      15 when "11101010011000",
                      15 when "11101010011001",
                      15 when "11101010011010",
                      15 when "11101010011011",
                      15 when "11101010011100",
                      15 when "11101010011101",
                      15 when "11101010011110",
                      15 when "11101010011111",
                      15 when "11101010100000",
                      15 when "11101010100001",
                      15 when "11101010100010",
                      15 when "11101010100011",
                      15 when "11101010100100",
                      15 when "11101010100101",
                      15 when "11101010100110",
                      15 when "11101010100111",
                      15 when "11101010101000",
                      15 when "11101010101001",
                      15 when "11101010101010",
                      15 when "11101010101011",
                      15 when "11101010101100",
                      15 when "11101010101101",
                      15 when "11101010101110",
                      15 when "11101010101111",
                      15 when "11101010110000",
                      15 when "11101010110001",
                      15 when "11101010110010",
                      15 when "11101010110011",
                      15 when "11101010110100",
                      15 when "11101010110101",
                      15 when "11101010110110",
                      15 when "11101010110111",
                      15 when "11101010111000",
                      15 when "11101010111001",
                      15 when "11101010111010",
                      15 when "11101010111011",
                      15 when "11101010111100",
                      15 when "11101010111101",
                      15 when "11101010111110",
                      15 when "11101010111111",
                      15 when "11101011000000",
                      15 when "11101011000001",
                      15 when "11101011000010",
                      15 when "11101011000011",
                      15 when "11101011000100",
                      15 when "11101011000101",
                      15 when "11101011000110",
                      15 when "11101011000111",
                      15 when "11101011001000",
                      15 when "11101011001001",
                      15 when "11101011001010",
                      15 when "11101011001011",
                      15 when "11101011001100",
                      15 when "11101011001101",
                      15 when "11101011001110",
                      15 when "11101011001111",
                      15 when "11101011010000",
                      15 when "11101011010001",
                      15 when "11101011010010",
                      15 when "11101011010011",
                      15 when "11101011010100",
                      15 when "11101011010101",
                      15 when "11101011010110",
                      15 when "11101011010111",
                      15 when "11101011011000",
                      15 when "11101011011001",
                      15 when "11101011011010",
                      15 when "11101011011011",
                      15 when "11101011011100",
                      15 when "11101011011101",
                      15 when "11101011011110",
                      15 when "11101011011111",
                      15 when "11101011100000",
                      15 when "11101011100001",
                      15 when "11101011100010",
                      15 when "11101011100011",
                      15 when "11101011100100",
                      15 when "11101011100101",
                      15 when "11101011100110",
                      15 when "11101011100111",
                      15 when "11101011101000",
                      15 when "11101011101001",
                      15 when "11101011101010",
                      15 when "11101011101011",
                      15 when "11101011101100",
                      15 when "11101011101101",
                      15 when "11101011101110",
                      15 when "11101011101111",
                      15 when "11101011110000",
                      15 when "11101011110001",
                      15 when "11101011110010",
                      15 when "11101011110011",
                      15 when "11101011110100",
                      15 when "11101011110101",
                      15 when "11101011110110",
                      15 when "11101011110111",
                      15 when "11101011111000",
                      15 when "11101011111001",
                      15 when "11101011111010",
                      15 when "11101011111011",
                      15 when "11101011111100",
                      15 when "11101011111101",
                      15 when "11101011111110",
                      15 when "11101011111111",
                      15 when "11101100000000",
                      15 when "11101100000001",
                      15 when "11101100000010",
                      15 when "11101100000011",
                      15 when "11101100000100",
                      15 when "11101100000101",
                      15 when "11101100000110",
                      15 when "11101100000111",
                      15 when "11101100001000",
                      15 when "11101100001001",
                      15 when "11101100001010",
                      15 when "11101100001011",
                      15 when "11101100001100",
                      15 when "11101100001101",
                      15 when "11101100001110",
                      15 when "11101100001111",
                      15 when "11101100010000",
                      15 when "11101100010001",
                      15 when "11101100010010",
                      15 when "11101100010011",
                      15 when "11101100010100",
                      15 when "11101100010101",
                      15 when "11101100010110",
                      15 when "11101100010111",
                      15 when "11101100011000",
                      15 when "11101100011001",
                      15 when "11101100011010",
                      15 when "11101100011011",
                      15 when "11101100011100",
                      15 when "11101100011101",
                      15 when "11101100011110",
                      15 when "11101100011111",
                      15 when "11101100100000",
                      15 when "11101100100001",
                      15 when "11101100100010",
                      15 when "11101100100011",
                      15 when "11101100100100",
                      15 when "11101100100101",
                      15 when "11101100100110",
                      15 when "11101100100111",
                      15 when "11101100101000",
                      15 when "11101100101001",
                      15 when "11101100101010",
                      15 when "11101100101011",
                      15 when "11101100101100",
                      15 when "11101100101101",
                      15 when "11101100101110",
                      15 when "11101100101111",
                      15 when "11101100110000",
                      15 when "11101100110001",
                      14 when "11101100110010",
                      14 when "11101100110011",
                      14 when "11101100110100",
                      14 when "11101100110101",
                      14 when "11101100110110",
                      14 when "11101100110111",
                      14 when "11101100111000",
                      14 when "11101100111001",
                      14 when "11101100111010",
                      14 when "11101100111011",
                      14 when "11101100111100",
                      14 when "11101100111101",
                      14 when "11101100111110",
                      14 when "11101100111111",
                      14 when "11101101000000",
                      14 when "11101101000001",
                      14 when "11101101000010",
                      14 when "11101101000011",
                      14 when "11101101000100",
                      14 when "11101101000101",
                      14 when "11101101000110",
                      14 when "11101101000111",
                      14 when "11101101001000",
                      14 when "11101101001001",
                      14 when "11101101001010",
                      14 when "11101101001011",
                      14 when "11101101001100",
                      14 when "11101101001101",
                      14 when "11101101001110",
                      14 when "11101101001111",
                      14 when "11101101010000",
                      14 when "11101101010001",
                      14 when "11101101010010",
                      14 when "11101101010011",
                      14 when "11101101010100",
                      14 when "11101101010101",
                      14 when "11101101010110",
                      14 when "11101101010111",
                      14 when "11101101011000",
                      14 when "11101101011001",
                      14 when "11101101011010",
                      14 when "11101101011011",
                      14 when "11101101011100",
                      14 when "11101101011101",
                      14 when "11101101011110",
                      14 when "11101101011111",
                      14 when "11101101100000",
                      14 when "11101101100001",
                      14 when "11101101100010",
                      14 when "11101101100011",
                      14 when "11101101100100",
                      14 when "11101101100101",
                      14 when "11101101100110",
                      14 when "11101101100111",
                      14 when "11101101101000",
                      14 when "11101101101001",
                      14 when "11101101101010",
                      14 when "11101101101011",
                      14 when "11101101101100",
                      14 when "11101101101101",
                      14 when "11101101101110",
                      14 when "11101101101111",
                      14 when "11101101110000",
                      14 when "11101101110001",
                      14 when "11101101110010",
                      14 when "11101101110011",
                      14 when "11101101110100",
                      14 when "11101101110101",
                      14 when "11101101110110",
                      14 when "11101101110111",
                      14 when "11101101111000",
                      14 when "11101101111001",
                      14 when "11101101111010",
                      14 when "11101101111011",
                      14 when "11101101111100",
                      14 when "11101101111101",
                      14 when "11101101111110",
                      14 when "11101101111111",
                      14 when "11101110000000",
                      14 when "11101110000001",
                      14 when "11101110000010",
                      14 when "11101110000011",
                      14 when "11101110000100",
                      14 when "11101110000101",
                      14 when "11101110000110",
                      14 when "11101110000111",
                      14 when "11101110001000",
                      14 when "11101110001001",
                      14 when "11101110001010",
                      14 when "11101110001011",
                      14 when "11101110001100",
                      14 when "11101110001101",
                      14 when "11101110001110",
                      14 when "11101110001111",
                      14 when "11101110010000",
                      14 when "11101110010001",
                      14 when "11101110010010",
                      14 when "11101110010011",
                      14 when "11101110010100",
                      14 when "11101110010101",
                      14 when "11101110010110",
                      14 when "11101110010111",
                      14 when "11101110011000",
                      14 when "11101110011001",
                      14 when "11101110011010",
                      14 when "11101110011011",
                      14 when "11101110011100",
                      14 when "11101110011101",
                      14 when "11101110011110",
                      14 when "11101110011111",
                      14 when "11101110100000",
                      14 when "11101110100001",
                      14 when "11101110100010",
                      14 when "11101110100011",
                      14 when "11101110100100",
                      14 when "11101110100101",
                      14 when "11101110100110",
                      14 when "11101110100111",
                      14 when "11101110101000",
                      14 when "11101110101001",
                      14 when "11101110101010",
                      14 when "11101110101011",
                      14 when "11101110101100",
                      14 when "11101110101101",
                      14 when "11101110101110",
                      14 when "11101110101111",
                      14 when "11101110110000",
                      14 when "11101110110001",
                      14 when "11101110110010",
                      14 when "11101110110011",
                      14 when "11101110110100",
                      14 when "11101110110101",
                      14 when "11101110110110",
                      14 when "11101110110111",
                      14 when "11101110111000",
                      14 when "11101110111001",
                      14 when "11101110111010",
                      14 when "11101110111011",
                      14 when "11101110111100",
                      14 when "11101110111101",
                      14 when "11101110111110",
                      14 when "11101110111111",
                      14 when "11101111000000",
                      14 when "11101111000001",
                      14 when "11101111000010",
                      14 when "11101111000011",
                      14 when "11101111000100",
                      14 when "11101111000101",
                      14 when "11101111000110",
                      14 when "11101111000111",
                      14 when "11101111001000",
                      14 when "11101111001001",
                      14 when "11101111001010",
                      14 when "11101111001011",
                      14 when "11101111001100",
                      14 when "11101111001101",
                      14 when "11101111001110",
                      14 when "11101111001111",
                      14 when "11101111010000",
                      14 when "11101111010001",
                      14 when "11101111010010",
                      14 when "11101111010011",
                      14 when "11101111010100",
                      14 when "11101111010101",
                      14 when "11101111010110",
                      14 when "11101111010111",
                      14 when "11101111011000",
                      14 when "11101111011001",
                      14 when "11101111011010",
                      14 when "11101111011011",
                      14 when "11101111011100",
                      14 when "11101111011101",
                      14 when "11101111011110",
                      14 when "11101111011111",
                      14 when "11101111100000",
                      14 when "11101111100001",
                      14 when "11101111100010",
                      14 when "11101111100011",
                      14 when "11101111100100",
                      14 when "11101111100101",
                      14 when "11101111100110",
                      14 when "11101111100111",
                      14 when "11101111101000",
                      14 when "11101111101001",
                      14 when "11101111101010",
                      14 when "11101111101011",
                      14 when "11101111101100",
                      14 when "11101111101101",
                      14 when "11101111101110",
                      14 when "11101111101111",
                      14 when "11101111110000",
                      14 when "11101111110001",
                      14 when "11101111110010",
                      14 when "11101111110011",
                      14 when "11101111110100",
                      14 when "11101111110101",
                      14 when "11101111110110",
                      14 when "11101111110111",
                      14 when "11101111111000",
                      14 when "11101111111001",
                      14 when "11101111111010",
                      14 when "11101111111011",
                      14 when "11101111111100",
                      14 when "11101111111101",
                      14 when "11101111111110",
                      14 when "11101111111111",
                      14 when "11110000000000",
                      14 when "11110000000001",
                      14 when "11110000000010",
                      14 when "11110000000011",
                      14 when "11110000000100",
                      14 when "11110000000101",
                      14 when "11110000000110",
                      14 when "11110000000111",
                      14 when "11110000001000",
                      14 when "11110000001001",
                      14 when "11110000001010",
                      14 when "11110000001011",
                      14 when "11110000001100",
                      14 when "11110000001101",
                      14 when "11110000001110",
                      14 when "11110000001111",
                      14 when "11110000010000",
                      14 when "11110000010001",
                      14 when "11110000010010",
                      14 when "11110000010011",
                      14 when "11110000010100",
                      14 when "11110000010101",
                      14 when "11110000010110",
                      14 when "11110000010111",
                      14 when "11110000011000",
                      14 when "11110000011001",
                      14 when "11110000011010",
                      14 when "11110000011011",
                      14 when "11110000011100",
                      14 when "11110000011101",
                      14 when "11110000011110",
                      14 when "11110000011111",
                      14 when "11110000100000",
                      14 when "11110000100001",
                      14 when "11110000100010",
                      14 when "11110000100011",
                      14 when "11110000100100",
                      14 when "11110000100101",
                      14 when "11110000100110",
                      14 when "11110000100111",
                      14 when "11110000101000",
                      14 when "11110000101001",
                      14 when "11110000101010",
                      14 when "11110000101011",
                      14 when "11110000101100",
                      14 when "11110000101101",
                      14 when "11110000101110",
                      14 when "11110000101111",
                      14 when "11110000110000",
                      14 when "11110000110001",
                      14 when "11110000110010",
                      14 when "11110000110011",
                      14 when "11110000110100",
                      14 when "11110000110101",
                      14 when "11110000110110",
                      14 when "11110000110111",
                      14 when "11110000111000",
                      14 when "11110000111001",
                      14 when "11110000111010",
                      14 when "11110000111011",
                      14 when "11110000111100",
                      14 when "11110000111101",
                      14 when "11110000111110",
                      14 when "11110000111111",
                      14 when "11110001000000",
                      14 when "11110001000001",
                      14 when "11110001000010",
                      14 when "11110001000011",
                      14 when "11110001000100",
                      14 when "11110001000101",
                      14 when "11110001000110",
                      14 when "11110001000111",
                      14 when "11110001001000",
                      14 when "11110001001001",
                      14 when "11110001001010",
                      14 when "11110001001011",
                      14 when "11110001001100",
                      14 when "11110001001101",
                      14 when "11110001001110",
                      14 when "11110001001111",
                      14 when "11110001010000",
                      14 when "11110001010001",
                      14 when "11110001010010",
                      14 when "11110001010011",
                      14 when "11110001010100",
                      14 when "11110001010101",
                      14 when "11110001010110",
                      14 when "11110001010111",
                      14 when "11110001011000",
                      14 when "11110001011001",
                      14 when "11110001011010",
                      14 when "11110001011011",
                      14 when "11110001011100",
                      14 when "11110001011101",
                      14 when "11110001011110",
                      14 when "11110001011111",
                      14 when "11110001100000",
                      14 when "11110001100001",
                      14 when "11110001100010",
                      14 when "11110001100011",
                      14 when "11110001100100",
                      14 when "11110001100101",
                      14 when "11110001100110",
                      14 when "11110001100111",
                      14 when "11110001101000",
                      14 when "11110001101001",
                      14 when "11110001101010",
                      14 when "11110001101011",
                      14 when "11110001101100",
                      14 when "11110001101101",
                      14 when "11110001101110",
                      14 when "11110001101111",
                      14 when "11110001110000",
                      14 when "11110001110001",
                      14 when "11110001110010",
                      14 when "11110001110011",
                      14 when "11110001110100",
                      14 when "11110001110101",
                      14 when "11110001110110",
                      14 when "11110001110111",
                      14 when "11110001111000",
                      14 when "11110001111001",
                      14 when "11110001111010",
                      14 when "11110001111011",
                      14 when "11110001111100",
                      14 when "11110001111101",
                      14 when "11110001111110",
                      14 when "11110001111111",
                      14 when "11110010000000",
                      14 when "11110010000001",
                      14 when "11110010000010",
                      14 when "11110010000011",
                      14 when "11110010000100",
                      14 when "11110010000101",
                      14 when "11110010000110",
                      14 when "11110010000111",
                      14 when "11110010001000",
                      14 when "11110010001001",
                      14 when "11110010001010",
                      14 when "11110010001011",
                      14 when "11110010001100",
                      14 when "11110010001101",
                      14 when "11110010001110",
                      14 when "11110010001111",
                      14 when "11110010010000",
                      14 when "11110010010001",
                      14 when "11110010010010",
                      14 when "11110010010011",
                      14 when "11110010010100",
                      14 when "11110010010101",
                      14 when "11110010010110",
                      14 when "11110010010111",
                      14 when "11110010011000",
                      14 when "11110010011001",
                      14 when "11110010011010",
                      14 when "11110010011011",
                      14 when "11110010011100",
                      14 when "11110010011101",
                      14 when "11110010011110",
                      14 when "11110010011111",
                      14 when "11110010100000",
                      14 when "11110010100001",
                      14 when "11110010100010",
                      14 when "11110010100011",
                      14 when "11110010100100",
                      14 when "11110010100101",
                      14 when "11110010100110",
                      14 when "11110010100111",
                      14 when "11110010101000",
                      14 when "11110010101001",
                      14 when "11110010101010",
                      14 when "11110010101011",
                      14 when "11110010101100",
                      14 when "11110010101101",
                      14 when "11110010101110",
                      14 when "11110010101111",
                      14 when "11110010110000",
                      14 when "11110010110001",
                      14 when "11110010110010",
                      14 when "11110010110011",
                      14 when "11110010110100",
                      14 when "11110010110101",
                      14 when "11110010110110",
                      14 when "11110010110111",
                      14 when "11110010111000",
                      14 when "11110010111001",
                      14 when "11110010111010",
                      14 when "11110010111011",
                      14 when "11110010111100",
                      14 when "11110010111101",
                      14 when "11110010111110",
                      14 when "11110010111111",
                      14 when "11110011000000",
                      14 when "11110011000001",
                      14 when "11110011000010",
                      14 when "11110011000011",
                      14 when "11110011000100",
                      14 when "11110011000101",
                      14 when "11110011000110",
                      14 when "11110011000111",
                      14 when "11110011001000",
                      14 when "11110011001001",
                      14 when "11110011001010",
                      14 when "11110011001011",
                      14 when "11110011001100",
                      14 when "11110011001101",
                      14 when "11110011001110",
                      14 when "11110011001111",
                      14 when "11110011010000",
                      14 when "11110011010001",
                      14 when "11110011010010",
                      14 when "11110011010011",
                      14 when "11110011010100",
                      14 when "11110011010101",
                      14 when "11110011010110",
                      14 when "11110011010111",
                      14 when "11110011011000",
                      14 when "11110011011001",
                      14 when "11110011011010",
                      14 when "11110011011011",
                      14 when "11110011011100",
                      14 when "11110011011101",
                      14 when "11110011011110",
                      14 when "11110011011111",
                      14 when "11110011100000",
                      14 when "11110011100001",
                      14 when "11110011100010",
                      14 when "11110011100011",
                      14 when "11110011100100",
                      14 when "11110011100101",
                      14 when "11110011100110",
                      14 when "11110011100111",
                      14 when "11110011101000",
                      14 when "11110011101001",
                      14 when "11110011101010",
                      14 when "11110011101011",
                      14 when "11110011101100",
                      14 when "11110011101101",
                      14 when "11110011101110",
                      14 when "11110011101111",
                      14 when "11110011110000",
                      14 when "11110011110001",
                      14 when "11110011110010",
                      14 when "11110011110011",
                      14 when "11110011110100",
                      14 when "11110011110101",
                      14 when "11110011110110",
                      14 when "11110011110111",
                      14 when "11110011111000",
                      14 when "11110011111001",
                      14 when "11110011111010",
                      14 when "11110011111011",
                      14 when "11110011111100",
                      14 when "11110011111101",
                      14 when "11110011111110",
                      14 when "11110011111111",
                      14 when "11110100000000",
                      14 when "11110100000001",
                      14 when "11110100000010",
                      14 when "11110100000011",
                      14 when "11110100000100",
                      14 when "11110100000101",
                      14 when "11110100000110",
                      14 when "11110100000111",
                      14 when "11110100001000",
                      14 when "11110100001001",
                      14 when "11110100001010",
                      14 when "11110100001011",
                      14 when "11110100001100",
                      14 when "11110100001101",
                      14 when "11110100001110",
                      14 when "11110100001111",
                      14 when "11110100010000",
                      14 when "11110100010001",
                      14 when "11110100010010",
                      14 when "11110100010011",
                      14 when "11110100010100",
                      14 when "11110100010101",
                      14 when "11110100010110",
                      14 when "11110100010111",
                      14 when "11110100011000",
                      14 when "11110100011001",
                      14 when "11110100011010",
                      14 when "11110100011011",
                      14 when "11110100011100",
                      14 when "11110100011101",
                      14 when "11110100011110",
                      14 when "11110100011111",
                      14 when "11110100100000",
                      14 when "11110100100001",
                      14 when "11110100100010",
                      14 when "11110100100011",
                      14 when "11110100100100",
                      14 when "11110100100101",
                      14 when "11110100100110",
                      14 when "11110100100111",
                      14 when "11110100101000",
                      14 when "11110100101001",
                      14 when "11110100101010",
                      14 when "11110100101011",
                      14 when "11110100101100",
                      14 when "11110100101101",
                      14 when "11110100101110",
                      14 when "11110100101111",
                      14 when "11110100110000",
                      14 when "11110100110001",
                      14 when "11110100110010",
                      14 when "11110100110011",
                      14 when "11110100110100",
                      14 when "11110100110101",
                      14 when "11110100110110",
                      14 when "11110100110111",
                      14 when "11110100111000",
                      14 when "11110100111001",
                      14 when "11110100111010",
                      14 when "11110100111011",
                      14 when "11110100111100",
                      14 when "11110100111101",
                      14 when "11110100111110",
                      14 when "11110100111111",
                      14 when "11110101000000",
                      14 when "11110101000001",
                      14 when "11110101000010",
                      14 when "11110101000011",
                      14 when "11110101000100",
                      14 when "11110101000101",
                      14 when "11110101000110",
                      14 when "11110101000111",
                      14 when "11110101001000",
                      14 when "11110101001001",
                      14 when "11110101001010",
                      14 when "11110101001011",
                      14 when "11110101001100",
                      14 when "11110101001101",
                      14 when "11110101001110",
                      14 when "11110101001111",
                      14 when "11110101010000",
                      14 when "11110101010001",
                      14 when "11110101010010",
                      14 when "11110101010011",
                      14 when "11110101010100",
                      14 when "11110101010101",
                      14 when "11110101010110",
                      14 when "11110101010111",
                      14 when "11110101011000",
                      14 when "11110101011001",
                      14 when "11110101011010",
                      14 when "11110101011011",
                      14 when "11110101011100",
                      14 when "11110101011101",
                      14 when "11110101011110",
                      14 when "11110101011111",
                      14 when "11110101100000",
                      14 when "11110101100001",
                      14 when "11110101100010",
                      14 when "11110101100011",
                      14 when "11110101100100",
                      14 when "11110101100101",
                      14 when "11110101100110",
                      14 when "11110101100111",
                      14 when "11110101101000",
                      14 when "11110101101001",
                      14 when "11110101101010",
                      14 when "11110101101011",
                      14 when "11110101101100",
                      14 when "11110101101101",
                      14 when "11110101101110",
                      14 when "11110101101111",
                      14 when "11110101110000",
                      14 when "11110101110001",
                      14 when "11110101110010",
                      14 when "11110101110011",
                      14 when "11110101110100",
                      14 when "11110101110101",
                      14 when "11110101110110",
                      14 when "11110101110111",
                      14 when "11110101111000",
                      14 when "11110101111001",
                      14 when "11110101111010",
                      14 when "11110101111011",
                      14 when "11110101111100",
                      14 when "11110101111101",
                      14 when "11110101111110",
                      14 when "11110101111111",
                      14 when "11110110000000",
                      14 when "11110110000001",
                      14 when "11110110000010",
                      14 when "11110110000011",
                      14 when "11110110000100",
                      14 when "11110110000101",
                      14 when "11110110000110",
                      14 when "11110110000111",
                      14 when "11110110001000",
                      14 when "11110110001001",
                      14 when "11110110001010",
                      14 when "11110110001011",
                      14 when "11110110001100",
                      14 when "11110110001101",
                      14 when "11110110001110",
                      14 when "11110110001111",
                      14 when "11110110010000",
                      14 when "11110110010001",
                      14 when "11110110010010",
                      14 when "11110110010011",
                      14 when "11110110010100",
                      14 when "11110110010101",
                      14 when "11110110010110",
                      14 when "11110110010111",
                      14 when "11110110011000",
                      14 when "11110110011001",
                      14 when "11110110011010",
                      14 when "11110110011011",
                      14 when "11110110011100",
                      14 when "11110110011101",
                      14 when "11110110011110",
                      14 when "11110110011111",
                      14 when "11110110100000",
                      14 when "11110110100001",
                      14 when "11110110100010",
                      14 when "11110110100011",
                      14 when "11110110100100",
                      14 when "11110110100101",
                      14 when "11110110100110",
                      14 when "11110110100111",
                      14 when "11110110101000",
                      14 when "11110110101001",
                      14 when "11110110101010",
                      14 when "11110110101011",
                      14 when "11110110101100",
                      14 when "11110110101101",
                      14 when "11110110101110",
                      14 when "11110110101111",
                      14 when "11110110110000",
                      14 when "11110110110001",
                      14 when "11110110110010",
                      14 when "11110110110011",
                      14 when "11110110110100",
                      14 when "11110110110101",
                      14 when "11110110110110",
                      14 when "11110110110111",
                      14 when "11110110111000",
                      14 when "11110110111001",
                      14 when "11110110111010",
                      14 when "11110110111011",
                      14 when "11110110111100",
                      14 when "11110110111101",
                      14 when "11110110111110",
                      14 when "11110110111111",
                      14 when "11110111000000",
                      14 when "11110111000001",
                      14 when "11110111000010",
                      14 when "11110111000011",
                      14 when "11110111000100",
                      14 when "11110111000101",
                      14 when "11110111000110",
                      14 when "11110111000111",
                      14 when "11110111001000",
                      14 when "11110111001001",
                      14 when "11110111001010",
                      14 when "11110111001011",
                      14 when "11110111001100",
                      14 when "11110111001101",
                      14 when "11110111001110",
                      14 when "11110111001111",
                      14 when "11110111010000",
                      14 when "11110111010001",
                      14 when "11110111010010",
                      14 when "11110111010011",
                      14 when "11110111010100",
                      14 when "11110111010101",
                      14 when "11110111010110",
                      14 when "11110111010111",
                      14 when "11110111011000",
                      14 when "11110111011001",
                      14 when "11110111011010",
                      14 when "11110111011011",
                      14 when "11110111011100",
                      14 when "11110111011101",
                      14 when "11110111011110",
                      14 when "11110111011111",
                      14 when "11110111100000",
                      14 when "11110111100001",
                      14 when "11110111100010",
                      14 when "11110111100011",
                      14 when "11110111100100",
                      14 when "11110111100101",
                      14 when "11110111100110",
                      14 when "11110111100111",
                      14 when "11110111101000",
                      14 when "11110111101001",
                      14 when "11110111101010",
                      14 when "11110111101011",
                      14 when "11110111101100",
                      14 when "11110111101101",
                      14 when "11110111101110",
                      14 when "11110111101111",
                      14 when "11110111110000",
                      14 when "11110111110001",
                      14 when "11110111110010",
                      14 when "11110111110011",
                      14 when "11110111110100",
                      14 when "11110111110101",
                      14 when "11110111110110",
                      14 when "11110111110111",
                      14 when "11110111111000",
                      14 when "11110111111001",
                      14 when "11110111111010",
                      14 when "11110111111011",
                      14 when "11110111111100",
                      14 when "11110111111101",
                      14 when "11110111111110",
                      14 when "11110111111111",
                      14 when "11111000000000",
                      14 when "11111000000001",
                      14 when "11111000000010",
                      14 when "11111000000011",
                      14 when "11111000000100",
                      14 when "11111000000101",
                      14 when "11111000000110",
                      14 when "11111000000111",
                      14 when "11111000001000",
                      14 when "11111000001001",
                      14 when "11111000001010",
                      14 when "11111000001011",
                      14 when "11111000001100",
                      14 when "11111000001101",
                      14 when "11111000001110",
                      14 when "11111000001111",
                      14 when "11111000010000",
                      14 when "11111000010001",
                      14 when "11111000010010",
                      14 when "11111000010011",
                      14 when "11111000010100",
                      14 when "11111000010101",
                      14 when "11111000010110",
                      14 when "11111000010111",
                      14 when "11111000011000",
                      14 when "11111000011001",
                      14 when "11111000011010",
                      14 when "11111000011011",
                      14 when "11111000011100",
                      14 when "11111000011101",
                      14 when "11111000011110",
                      14 when "11111000011111",
                      14 when "11111000100000",
                      14 when "11111000100001",
                      14 when "11111000100010",
                      14 when "11111000100011",
                      14 when "11111000100100",
                      14 when "11111000100101",
                      14 when "11111000100110",
                      14 when "11111000100111",
                      14 when "11111000101000",
                      14 when "11111000101001",
                      14 when "11111000101010",
                      14 when "11111000101011",
                      14 when "11111000101100",
                      14 when "11111000101101",
                      14 when "11111000101110",
                      14 when "11111000101111",
                      14 when "11111000110000",
                      14 when "11111000110001",
                      14 when "11111000110010",
                      14 when "11111000110011",
                      14 when "11111000110100",
                      14 when "11111000110101",
                      14 when "11111000110110",
                      14 when "11111000110111",
                      14 when "11111000111000",
                      14 when "11111000111001",
                      14 when "11111000111010",
                      14 when "11111000111011",
                      14 when "11111000111100",
                      14 when "11111000111101",
                      14 when "11111000111110",
                      14 when "11111000111111",
                      14 when "11111001000000",
                      14 when "11111001000001",
                      14 when "11111001000010",
                      14 when "11111001000011",
                      14 when "11111001000100",
                      14 when "11111001000101",
                      14 when "11111001000110",
                      14 when "11111001000111",
                      14 when "11111001001000",
                      14 when "11111001001001",
                      14 when "11111001001010",
                      14 when "11111001001011",
                      14 when "11111001001100",
                      14 when "11111001001101",
                      14 when "11111001001110",
                      14 when "11111001001111",
                      14 when "11111001010000",
                      14 when "11111001010001",
                      14 when "11111001010010",
                      14 when "11111001010011",
                      14 when "11111001010100",
                      14 when "11111001010101",
                      14 when "11111001010110",
                      14 when "11111001010111",
                      14 when "11111001011000",
                      14 when "11111001011001",
                      14 when "11111001011010",
                      14 when "11111001011011",
                      14 when "11111001011100",
                      14 when "11111001011101",
                      14 when "11111001011110",
                      14 when "11111001011111",
                      14 when "11111001100000",
                      14 when "11111001100001",
                      14 when "11111001100010",
                      14 when "11111001100011",
                      14 when "11111001100100",
                      14 when "11111001100101",
                      14 when "11111001100110",
                      14 when "11111001100111",
                      14 when "11111001101000",
                      14 when "11111001101001",
                      14 when "11111001101010",
                      14 when "11111001101011",
                      14 when "11111001101100",
                      14 when "11111001101101",
                      14 when "11111001101110",
                      14 when "11111001101111",
                      14 when "11111001110000",
                      14 when "11111001110001",
                      14 when "11111001110010",
                      14 when "11111001110011",
                      14 when "11111001110100",
                      14 when "11111001110101",
                      14 when "11111001110110",
                      14 when "11111001110111",
                      14 when "11111001111000",
                      14 when "11111001111001",
                      14 when "11111001111010",
                      14 when "11111001111011",
                      14 when "11111001111100",
                      14 when "11111001111101",
                      14 when "11111001111110",
                      14 when "11111001111111",
                      14 when "11111010000000",
                      14 when "11111010000001",
                      14 when "11111010000010",
                      14 when "11111010000011",
                      14 when "11111010000100",
                      14 when "11111010000101",
                      14 when "11111010000110",
                      14 when "11111010000111",
                      14 when "11111010001000",
                      14 when "11111010001001",
                      14 when "11111010001010",
                      14 when "11111010001011",
                      14 when "11111010001100",
                      14 when "11111010001101",
                      14 when "11111010001110",
                      14 when "11111010001111",
                      14 when "11111010010000",
                      14 when "11111010010001",
                      14 when "11111010010010",
                      14 when "11111010010011",
                      14 when "11111010010100",
                      14 when "11111010010101",
                      14 when "11111010010110",
                      14 when "11111010010111",
                      14 when "11111010011000",
                      14 when "11111010011001",
                      14 when "11111010011010",
                      14 when "11111010011011",
                      14 when "11111010011100",
                      14 when "11111010011101",
                      14 when "11111010011110",
                      14 when "11111010011111",
                      14 when "11111010100000",
                      14 when "11111010100001",
                      14 when "11111010100010",
                      14 when "11111010100011",
                      14 when "11111010100100",
                      14 when "11111010100101",
                      14 when "11111010100110",
                      14 when "11111010100111",
                      14 when "11111010101000",
                      14 when "11111010101001",
                      14 when "11111010101010",
                      14 when "11111010101011",
                      14 when "11111010101100",
                      14 when "11111010101101",
                      14 when "11111010101110",
                      14 when "11111010101111",
                      14 when "11111010110000",
                      14 when "11111010110001",
                      14 when "11111010110010",
                      14 when "11111010110011",
                      14 when "11111010110100",
                      14 when "11111010110101",
                      14 when "11111010110110",
                      14 when "11111010110111",
                      14 when "11111010111000",
                      14 when "11111010111001",
                      14 when "11111010111010",
                      14 when "11111010111011",
                      14 when "11111010111100",
                      14 when "11111010111101",
                      14 when "11111010111110",
                      14 when "11111010111111",
                      14 when "11111011000000",
                      14 when "11111011000001",
                      14 when "11111011000010",
                      14 when "11111011000011",
                      14 when "11111011000100",
                      14 when "11111011000101",
                      14 when "11111011000110",
                      14 when "11111011000111",
                      14 when "11111011001000",
                      14 when "11111011001001",
                      14 when "11111011001010",
                      14 when "11111011001011",
                      14 when "11111011001100",
                      14 when "11111011001101",
                      14 when "11111011001110",
                      14 when "11111011001111",
                      14 when "11111011010000",
                      14 when "11111011010001",
                      14 when "11111011010010",
                      14 when "11111011010011",
                      14 when "11111011010100",
                      14 when "11111011010101",
                      14 when "11111011010110",
                      14 when "11111011010111",
                      14 when "11111011011000",
                      14 when "11111011011001",
                      14 when "11111011011010",
                      14 when "11111011011011",
                      14 when "11111011011100",
                      14 when "11111011011101",
                      14 when "11111011011110",
                      14 when "11111011011111",
                      14 when "11111011100000",
                      14 when "11111011100001",
                      14 when "11111011100010",
                      14 when "11111011100011",
                      14 when "11111011100100",
                      14 when "11111011100101",
                      14 when "11111011100110",
                      14 when "11111011100111",
                      14 when "11111011101000",
                      14 when "11111011101001",
                      14 when "11111011101010",
                      14 when "11111011101011",
                      14 when "11111011101100",
                      14 when "11111011101101",
                      14 when "11111011101110",
                      14 when "11111011101111",
                      14 when "11111011110000",
                      14 when "11111011110001",
                      14 when "11111011110010",
                      14 when "11111011110011",
                      14 when "11111011110100",
                      14 when "11111011110101",
                      14 when "11111011110110",
                      14 when "11111011110111",
                      14 when "11111011111000",
                      14 when "11111011111001",
                      14 when "11111011111010",
                      14 when "11111011111011",
                      14 when "11111011111100",
                      14 when "11111011111101",
                      14 when "11111011111110",
                      14 when "11111011111111",
                      14 when "11111100000000",
                      14 when "11111100000001",
                      14 when "11111100000010",
                      14 when "11111100000011",
                      14 when "11111100000100",
                      14 when "11111100000101",
                      14 when "11111100000110",
                      14 when "11111100000111",
                      14 when "11111100001000",
                      14 when "11111100001001",
                      14 when "11111100001010",
                      14 when "11111100001011",
                      14 when "11111100001100",
                      14 when "11111100001101",
                      14 when "11111100001110",
                      14 when "11111100001111",
                      14 when "11111100010000",
                      14 when "11111100010001",
                      14 when "11111100010010",
                      14 when "11111100010011",
                      14 when "11111100010100",
                      14 when "11111100010101",
                      14 when "11111100010110",
                      14 when "11111100010111",
                      14 when "11111100011000",
                      14 when "11111100011001",
                      14 when "11111100011010",
                      14 when "11111100011011",
                      14 when "11111100011100",
                      14 when "11111100011101",
                      14 when "11111100011110",
                      14 when "11111100011111",
                      14 when "11111100100000",
                      14 when "11111100100001",
                      14 when "11111100100010",
                      14 when "11111100100011",
                      14 when "11111100100100",
                      14 when "11111100100101",
                      14 when "11111100100110",
                      14 when "11111100100111",
                      14 when "11111100101000",
                      14 when "11111100101001",
                      14 when "11111100101010",
                      14 when "11111100101011",
                      14 when "11111100101100",
                      14 when "11111100101101",
                      14 when "11111100101110",
                      14 when "11111100101111",
                      14 when "11111100110000",
                      14 when "11111100110001",
                      14 when "11111100110010",
                      14 when "11111100110011",
                      14 when "11111100110100",
                      14 when "11111100110101",
                      14 when "11111100110110",
                      14 when "11111100110111",
                      14 when "11111100111000",
                      14 when "11111100111001",
                      14 when "11111100111010",
                      14 when "11111100111011",
                      14 when "11111100111100",
                      14 when "11111100111101",
                      14 when "11111100111110",
                      14 when "11111100111111",
                      14 when "11111101000000",
                      14 when "11111101000001",
                      14 when "11111101000010",
                      14 when "11111101000011",
                      14 when "11111101000100",
                      14 when "11111101000101",
                      14 when "11111101000110",
                      14 when "11111101000111",
                      14 when "11111101001000",
                      14 when "11111101001001",
                      14 when "11111101001010",
                      14 when "11111101001011",
                      14 when "11111101001100",
                      14 when "11111101001101",
                      14 when "11111101001110",
                      14 when "11111101001111",
                      14 when "11111101010000",
                      14 when "11111101010001",
                      14 when "11111101010010",
                      14 when "11111101010011",
                      14 when "11111101010100",
                      14 when "11111101010101",
                      14 when "11111101010110",
                      14 when "11111101010111",
                      14 when "11111101011000",
                      14 when "11111101011001",
                      14 when "11111101011010",
                      14 when "11111101011011",
                      14 when "11111101011100",
                      14 when "11111101011101",
                      14 when "11111101011110",
                      14 when "11111101011111",
                      14 when "11111101100000",
                      14 when "11111101100001",
                      14 when "11111101100010",
                      14 when "11111101100011",
                      14 when "11111101100100",
                      14 when "11111101100101",
                      14 when "11111101100110",
                      14 when "11111101100111",
                      14 when "11111101101000",
                      14 when "11111101101001",
                      14 when "11111101101010",
                      14 when "11111101101011",
                      14 when "11111101101100",
                      14 when "11111101101101",
                      14 when "11111101101110",
                      14 when "11111101101111",
                      14 when "11111101110000",
                      14 when "11111101110001",
                      14 when "11111101110010",
                      14 when "11111101110011",
                      14 when "11111101110100",
                      14 when "11111101110101",
                      14 when "11111101110110",
                      14 when "11111101110111",
                      14 when "11111101111000",
                      14 when "11111101111001",
                      14 when "11111101111010",
                      14 when "11111101111011",
                      14 when "11111101111100",
                      14 when "11111101111101",
                      14 when "11111101111110",
                      14 when "11111101111111",
                      14 when "11111110000000",
                      14 when "11111110000001",
                      14 when "11111110000010",
                      14 when "11111110000011",
                      14 when "11111110000100",
                      14 when "11111110000101",
                      14 when "11111110000110",
                      14 when "11111110000111",
                      14 when "11111110001000",
                      14 when "11111110001001",
                      14 when "11111110001010",
                      14 when "11111110001011",
                      14 when "11111110001100",
                      14 when "11111110001101",
                      14 when "11111110001110",
                      14 when "11111110001111",
                      14 when "11111110010000",
                      14 when "11111110010001",
                      14 when "11111110010010",
                      14 when "11111110010011",
                      14 when "11111110010100",
                      13 when "11111110010101",
                      13 when "11111110010110",
                      13 when "11111110010111",
                      13 when "11111110011000",
                      13 when "11111110011001",
                      13 when "11111110011010",
                      13 when "11111110011011",
                      13 when "11111110011100",
                      13 when "11111110011101",
                      13 when "11111110011110",
                      13 when "11111110011111",
                      13 when "11111110100000",
                      13 when "11111110100001",
                      13 when "11111110100010",
                      13 when "11111110100011",
                      13 when "11111110100100",
                      13 when "11111110100101",
                      13 when "11111110100110",
                      13 when "11111110100111",
                      13 when "11111110101000",
                      13 when "11111110101001",
                      13 when "11111110101010",
                      13 when "11111110101011",
                      13 when "11111110101100",
                      13 when "11111110101101",
                      13 when "11111110101110",
                      13 when "11111110101111",
                      13 when "11111110110000",
                      13 when "11111110110001",
                      13 when "11111110110010",
                      13 when "11111110110011",
                      13 when "11111110110100",
                      13 when "11111110110101",
                      13 when "11111110110110",
                      13 when "11111110110111",
                      13 when "11111110111000",
                      13 when "11111110111001",
                      13 when "11111110111010",
                      13 when "11111110111011",
                      13 when "11111110111100",
                      13 when "11111110111101",
                      13 when "11111110111110",
                      13 when "11111110111111",
                      13 when "11111111000000",
                      13 when "11111111000001",
                      13 when "11111111000010",
                      13 when "11111111000011",
                      13 when "11111111000100",
                      13 when "11111111000101",
                      13 when "11111111000110",
                      13 when "11111111000111",
                      13 when "11111111001000",
                      13 when "11111111001001",
                      13 when "11111111001010",
                      13 when "11111111001011",
                      13 when "11111111001100",
                      13 when "11111111001101",
                      13 when "11111111001110",
                      13 when "11111111001111",
                      13 when "11111111010000",
                      13 when "11111111010001",
                      13 when "11111111010010",
                      13 when "11111111010011",
                      13 when "11111111010100",
                      13 when "11111111010101",
                      13 when "11111111010110",
                      13 when "11111111010111",
                      13 when "11111111011000",
                      13 when "11111111011001",
                      13 when "11111111011010",
                      13 when "11111111011011",
                      13 when "11111111011100",
                      13 when "11111111011101",
                      13 when "11111111011110",
                      13 when "11111111011111",
                      13 when "11111111100000",
                      13 when "11111111100001",
                      13 when "11111111100010",
                      13 when "11111111100011",
                      13 when "11111111100100",
                      13 when "11111111100101",
                      13 when "11111111100110",
                      13 when "11111111100111",
                      13 when "11111111101000",
                      13 when "11111111101001",
                      13 when "11111111101010",
                      13 when "11111111101011",
                      13 when "11111111101100",
                      13 when "11111111101101",
                      13 when "11111111101110",
                      13 when "11111111101111",
                      13 when "11111111110000",
                      13 when "11111111110001",
                      13 when "11111111110010",
                      13 when "11111111110011",
                      13 when "11111111110100",
                      13 when "11111111110101",
                      13 when "11111111110110",
                      13 when "11111111110111",
                      13 when "11111111111000",
                      13 when "11111111111001",
                      13 when "11111111111010",
                      13 when "11111111111011",
                      13 when "11111111111100",
                      13 when "11111111111101",
                      13 when "11111111111110",
                      13 when "11111111111111",
                      0 when others;

end Behavioral;
