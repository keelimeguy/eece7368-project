-- Keelin Becker-Wheeler
-- lut_note_freq.vhd

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;

entity lut_note_freq is
    port (
        note_value : in  std_logic_vector(7 downto 0);
        freq_value : out std_logic_vector(13 downto 0)
    );
end lut_note_freq;

architecture Behavioral of lut_note_freq is
begin
    with note_value select
        freq_value <= "00000000001000" when "00000000",
                      "00000000001001" when "00000001",
                      "00000000001001" when "00000010",
                      "00000000001010" when "00000011",
                      "00000000001010" when "00000100",
                      "00000000001011" when "00000101",
                      "00000000001100" when "00000110",
                      "00000000001100" when "00000111",
                      "00000000001101" when "00001000",
                      "00000000001110" when "00001001",
                      "00000000001111" when "00001010",
                      "00000000001111" when "00001011",
                      "00000000010000" when "00001100",
                      "00000000010001" when "00001101",
                      "00000000010010" when "00001110",
                      "00000000010011" when "00001111",
                      "00000000010101" when "00010000",
                      "00000000010110" when "00010001",
                      "00000000010111" when "00010010",
                      "00000000011001" when "00010011",
                      "00000000011010" when "00010100",
                      "00000000011100" when "00010101",
                      "00000000011101" when "00010110",
                      "00000000011111" when "00010111",
                      "00000000100001" when "00011000",
                      "00000000100011" when "00011001",
                      "00000000100101" when "00011010",
                      "00000000100111" when "00011011",
                      "00000000101001" when "00011100",
                      "00000000101100" when "00011101",
                      "00000000101110" when "00011110",
                      "00000000110001" when "00011111",
                      "00000000110100" when "00100000",
                      "00000000110111" when "00100001",
                      "00000000111010" when "00100010",
                      "00000000111110" when "00100011",
                      "00000001000001" when "00100100",
                      "00000001000101" when "00100101",
                      "00000001001001" when "00100110",
                      "00000001001110" when "00100111",
                      "00000001010010" when "00101000",
                      "00000001010111" when "00101001",
                      "00000001011101" when "00101010",
                      "00000001100010" when "00101011",
                      "00000001101000" when "00101100",
                      "00000001101110" when "00101101",
                      "00000001110110" when "00101110",
                      "00000001111011" when "00101111",
                      "00000010000011" when "00110000",
                      "00000010001011" when "00110001",
                      "00000010010011" when "00110010",
                      "00000010011100" when "00110011",
                      "00000010100101" when "00110100",
                      "00000010101111" when "00110101",
                      "00000010111001" when "00110110",
                      "00000011000100" when "00110111",
                      "00000011010000" when "00111000",
                      "00000011011100" when "00111001",
                      "00000011101001" when "00111010",
                      "00000011110111" when "00111011",
                      "00000100000110" when "00111100",
                      "00000100010101" when "00111101",
                      "00000100100110" when "00111110",
                      "00000100110111" when "00111111",
                      "00000101001010" when "01000000",
                      "00000101011101" when "01000001",
                      "00000101110010" when "01000010",
                      "00000110001000" when "01000011",
                      "00000110011111" when "01000100",
                      "00000110111000" when "01000101",
                      "00000111010010" when "01000110",
                      "00000111101110" when "01000111",
                      "00001000001011" when "01001000",
                      "00001000101010" when "01001001",
                      "00001001001011" when "01001010",
                      "00001001101110" when "01001011",
                      "00001010010011" when "01001100",
                      "00001010111010" when "01001101",
                      "00001011100100" when "01001110",
                      "00001100010000" when "01001111",
                      "00001100111111" when "01010000",
                      "00001101110000" when "01010001",
                      "00001110100100" when "01010010",
                      "00001111011100" when "01010011",
                      "00010000010111" when "01010100",
                      "00010001010101" when "01010101",
                      "00010010010111" when "01010110",
                      "00010011011101" when "01010111",
                      "00010100100111" when "01011000",
                      "00010101110101" when "01011001",
                      "00010111001000" when "01011010",
                      "00011000100000" when "01011011",
                      "00011001111101" when "01011100",
                      "00011011100000" when "01011101",
                      "00011101001001" when "01011110",
                      "00011110111000" when "01011111",
                      "00100000101101" when "01100000",
                      "00100010101001" when "01100001",
                      "00100100101101" when "01100010",
                      "00100110111001" when "01100011",
                      "00101001001101" when "01100100",
                      "00101011101010" when "01100101",
                      "00101110010000" when "01100110",
                      "00110001000000" when "01100111",
                      "00110011111010" when "01101000",
                      "00110111000000" when "01101001",
                      "00111010010001" when "01101010",
                      "00111101101111" when "01101011",
                      "01000001011010" when "01101100",
                      "01000101010011" when "01101101",
                      "01001001011011" when "01101110",
                      "01001101110010" when "01101111",
                      "01010010011010" when "01110000",
                      "01010111010100" when "01110001",
                      "01011100100000" when "01110010",
                      "01100010000000" when "01110011",
                      "01100111110101" when "01110100",
                      "01101110000000" when "01110101",
                      "01110100100100" when "01110110",
                      "01111011011110" when "01110111",
                      "10000010110100" when "01111000",
                      "10001010100110" when "01111001",
                      "10010010110101" when "01111010",
                      "10011011100100" when "01111011",
                      "10100100110100" when "01111100",
                      "10101110100111" when "01111101",
                      "10111001000000" when "01111110",
                      "11000100000000" when "01111111",
                      "00000000000000" when others;
end Behavioral;
